

module test
(

);

  reg CLK;
  reg RESETN;
  wire irq;
  wire [32-1:0] maxi_awaddr;
  wire [8-1:0] maxi_awlen;
  wire [3-1:0] maxi_awsize;
  wire [2-1:0] maxi_awburst;
  wire [1-1:0] maxi_awlock;
  wire [4-1:0] maxi_awcache;
  wire [3-1:0] maxi_awprot;
  wire [4-1:0] maxi_awqos;
  wire [2-1:0] maxi_awuser;
  wire maxi_awvalid;
  reg maxi_awready;
  wire [32-1:0] maxi_wdata;
  wire [4-1:0] maxi_wstrb;
  wire maxi_wlast;
  wire maxi_wvalid;
  reg maxi_wready;
  reg [2-1:0] maxi_bresp;
  reg maxi_bvalid;
  wire maxi_bready;
  wire [32-1:0] maxi_araddr;
  wire [8-1:0] maxi_arlen;
  wire [3-1:0] maxi_arsize;
  wire [2-1:0] maxi_arburst;
  wire [1-1:0] maxi_arlock;
  wire [4-1:0] maxi_arcache;
  wire [3-1:0] maxi_arprot;
  wire [4-1:0] maxi_arqos;
  wire [2-1:0] maxi_aruser;
  wire maxi_arvalid;
  reg maxi_arready;
  reg [32-1:0] maxi_rdata;
  reg [2-1:0] maxi_rresp;
  reg maxi_rlast;
  reg maxi_rvalid;
  wire maxi_rready;
  reg [32-1:0] saxi_awaddr;
  reg [4-1:0] saxi_awcache;
  reg [3-1:0] saxi_awprot;
  reg saxi_awvalid;
  wire saxi_awready;
  reg [32-1:0] saxi_wdata;
  reg [4-1:0] saxi_wstrb;
  reg saxi_wvalid;
  wire saxi_wready;
  wire [2-1:0] saxi_bresp;
  wire saxi_bvalid;
  reg saxi_bready;
  reg [32-1:0] saxi_araddr;
  reg [4-1:0] saxi_arcache;
  reg [3-1:0] saxi_arprot;
  reg saxi_arvalid;
  wire saxi_arready;
  wire [32-1:0] saxi_rdata;
  wire [2-1:0] saxi_rresp;
  wire saxi_rvalid;
  reg saxi_rready;
  wire RST;
  assign RST = !RESETN;
  wire [32-1:0] memory_awaddr;
  wire [8-1:0] memory_awlen;
  wire [3-1:0] memory_awsize;
  wire [2-1:0] memory_awburst;
  wire [1-1:0] memory_awlock;
  wire [4-1:0] memory_awcache;
  wire [3-1:0] memory_awprot;
  wire [4-1:0] memory_awqos;
  wire [2-1:0] memory_awuser;
  wire memory_awvalid;
  reg memory_awready;
  wire [32-1:0] memory_wdata;
  wire [4-1:0] memory_wstrb;
  wire memory_wlast;
  wire memory_wvalid;
  wire memory_wready;
  wire [2-1:0] memory_bresp;
  reg memory_bvalid;
  wire memory_bready;
  assign memory_bresp = 0;
  wire [32-1:0] memory_araddr;
  wire [8-1:0] memory_arlen;
  wire [3-1:0] memory_arsize;
  wire [2-1:0] memory_arburst;
  wire [1-1:0] memory_arlock;
  wire [4-1:0] memory_arcache;
  wire [3-1:0] memory_arprot;
  wire [4-1:0] memory_arqos;
  wire [2-1:0] memory_aruser;
  wire memory_arvalid;
  reg memory_arready;
  reg [32-1:0] memory_rdata;
  wire [2-1:0] memory_rresp;
  reg memory_rlast;
  reg memory_rvalid;
  wire memory_rready;
  assign memory_rresp = 0;
  reg [32-1:0] _memory_waddr_fsm;
  localparam _memory_waddr_fsm_init = 0;
  reg [32-1:0] _memory_wdata_fsm;
  localparam _memory_wdata_fsm_init = 0;
  reg [32-1:0] _memory_raddr_fsm;
  localparam _memory_raddr_fsm_init = 0;
  reg [32-1:0] _memory_rdata_fsm;
  localparam _memory_rdata_fsm_init = 0;
  wire _memory_wreq_fifo_enq;
  wire [41-1:0] _memory_wreq_fifo_wdata;
  wire _memory_wreq_fifo_full;
  wire _memory_wreq_fifo_almost_full;
  wire _memory_wreq_fifo_deq;
  wire [41-1:0] _memory_wreq_fifo_rdata;
  wire _memory_wreq_fifo_empty;
  wire _memory_wreq_fifo_almost_empty;

  _memory_wreq_fifo
  inst__memory_wreq_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._memory_wreq_fifo_enq(_memory_wreq_fifo_enq),
    ._memory_wreq_fifo_wdata(_memory_wreq_fifo_wdata),
    ._memory_wreq_fifo_full(_memory_wreq_fifo_full),
    ._memory_wreq_fifo_almost_full(_memory_wreq_fifo_almost_full),
    ._memory_wreq_fifo_deq(_memory_wreq_fifo_deq),
    ._memory_wreq_fifo_rdata(_memory_wreq_fifo_rdata),
    ._memory_wreq_fifo_empty(_memory_wreq_fifo_empty),
    ._memory_wreq_fifo_almost_empty(_memory_wreq_fifo_almost_empty)
  );

  reg [4-1:0] count__memory_wreq_fifo;
  wire _memory_rreq_fifo_enq;
  wire [41-1:0] _memory_rreq_fifo_wdata;
  wire _memory_rreq_fifo_full;
  wire _memory_rreq_fifo_almost_full;
  wire _memory_rreq_fifo_deq;
  wire [41-1:0] _memory_rreq_fifo_rdata;
  wire _memory_rreq_fifo_empty;
  wire _memory_rreq_fifo_almost_empty;

  _memory_rreq_fifo
  inst__memory_rreq_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._memory_rreq_fifo_enq(_memory_rreq_fifo_enq),
    ._memory_rreq_fifo_wdata(_memory_rreq_fifo_wdata),
    ._memory_rreq_fifo_full(_memory_rreq_fifo_full),
    ._memory_rreq_fifo_almost_full(_memory_rreq_fifo_almost_full),
    ._memory_rreq_fifo_deq(_memory_rreq_fifo_deq),
    ._memory_rreq_fifo_rdata(_memory_rreq_fifo_rdata),
    ._memory_rreq_fifo_empty(_memory_rreq_fifo_empty),
    ._memory_rreq_fifo_almost_empty(_memory_rreq_fifo_almost_empty)
  );

  reg [4-1:0] count__memory_rreq_fifo;
  wire _memory_wdata_fifo_enq;
  wire [37-1:0] _memory_wdata_fifo_wdata;
  wire _memory_wdata_fifo_full;
  wire _memory_wdata_fifo_almost_full;
  wire _memory_wdata_fifo_deq;
  wire [37-1:0] _memory_wdata_fifo_rdata;
  wire _memory_wdata_fifo_empty;
  wire _memory_wdata_fifo_almost_empty;

  _memory_wdata_fifo
  inst__memory_wdata_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._memory_wdata_fifo_enq(_memory_wdata_fifo_enq),
    ._memory_wdata_fifo_wdata(_memory_wdata_fifo_wdata),
    ._memory_wdata_fifo_full(_memory_wdata_fifo_full),
    ._memory_wdata_fifo_almost_full(_memory_wdata_fifo_almost_full),
    ._memory_wdata_fifo_deq(_memory_wdata_fifo_deq),
    ._memory_wdata_fifo_rdata(_memory_wdata_fifo_rdata),
    ._memory_wdata_fifo_empty(_memory_wdata_fifo_empty),
    ._memory_wdata_fifo_almost_empty(_memory_wdata_fifo_almost_empty)
  );

  reg [4-1:0] count__memory_wdata_fifo;
  assign memory_wready = !_memory_wdata_fifo_almost_full;
  wire [32-1:0] pack_write_data_wdata_0;
  wire [4-1:0] pack_write_data_wstrb_1;
  wire [1-1:0] pack_write_data_wlast_2;
  assign pack_write_data_wdata_0 = memory_wdata;
  assign pack_write_data_wstrb_1 = memory_wstrb;
  assign pack_write_data_wlast_2 = memory_wlast;
  wire [37-1:0] pack_write_data_packed_3;
  assign pack_write_data_packed_3 = { pack_write_data_wlast_2, pack_write_data_wstrb_1, pack_write_data_wdata_0 };
  assign _memory_wdata_fifo_wdata = (memory_wvalid && memory_wready)? pack_write_data_packed_3 : 'hx;
  assign _memory_wdata_fifo_enq = (memory_wvalid && memory_wready)? memory_wvalid && memory_wready && !_memory_wdata_fifo_almost_full : 0;
  localparam _tmp_4 = 1;
  wire [_tmp_4-1:0] _tmp_5;
  assign _tmp_5 = !_memory_wdata_fifo_almost_full;
  reg [_tmp_4-1:0] __tmp_5_1;
  reg [8-1:0] _memory_mem [0:2**25-1];

  initial begin
    $readmemh("memimg_hello_nngen.out", _memory_mem);
  end

  reg [33-1:0] _write_count;
  reg [32-1:0] _write_addr;
  reg [33-1:0] _read_count;
  reg [32-1:0] _read_addr;
  reg [33-1:0] _sleep_interval_count;
  reg [33-1:0] _keep_sleep_count;
  wire [32-1:0] pack_write_req_global_addr_6;
  wire [9-1:0] pack_write_req_size_7;
  assign pack_write_req_global_addr_6 = memory_awaddr;
  assign pack_write_req_size_7 = memory_awlen + 1;
  wire [41-1:0] pack_write_req_packed_8;
  assign pack_write_req_packed_8 = { pack_write_req_global_addr_6, pack_write_req_size_7 };
  assign _memory_wreq_fifo_wdata = ((_memory_waddr_fsm == 11) && memory_awvalid && memory_awready)? pack_write_req_packed_8 : 'hx;
  assign _memory_wreq_fifo_enq = ((_memory_waddr_fsm == 11) && memory_awvalid && memory_awready)? (_memory_waddr_fsm == 11) && memory_awvalid && memory_awready && !_memory_wreq_fifo_almost_full : 0;
  localparam _tmp_9 = 1;
  wire [_tmp_9-1:0] _tmp_10;
  assign _tmp_10 = !_memory_wreq_fifo_almost_full;
  reg [_tmp_9-1:0] __tmp_10_1;
  wire [32-1:0] unpack_write_req_global_addr_11;
  wire [9-1:0] unpack_write_req_size_12;
  assign unpack_write_req_global_addr_11 = _memory_wreq_fifo_rdata[40:9];
  assign unpack_write_req_size_12 = _memory_wreq_fifo_rdata[8:0];
  assign _memory_wreq_fifo_deq = ((_memory_wdata_fsm == 0) && !_memory_wreq_fifo_empty && !_memory_wreq_fifo_empty)? 1 : 0;
  wire [32-1:0] pack_write_data_wdata_13;
  wire [4-1:0] pack_write_data_wstrb_14;
  wire [1-1:0] pack_write_data_wlast_15;
  assign pack_write_data_wdata_13 = _memory_wdata_fifo_rdata[31:0];
  assign pack_write_data_wstrb_14 = _memory_wdata_fifo_rdata[35:32];
  assign pack_write_data_wlast_15 = _memory_wdata_fifo_rdata[36];
  wire write_data_wvalid_16;
  assign write_data_wvalid_16 = !_memory_wdata_fifo_empty;
  wire write_data_wready_17;
  assign write_data_wready_17 = (_memory_wdata_fsm == 1) && (_sleep_interval_count != 15);
  assign _memory_wdata_fifo_deq = (write_data_wready_17 && !_memory_wdata_fifo_empty && !_memory_wdata_fifo_empty)? 1 : 0;
  wire [32-1:0] pack_read_req_global_addr_18;
  wire [9-1:0] pack_read_req_size_19;
  assign pack_read_req_global_addr_18 = memory_araddr;
  assign pack_read_req_size_19 = memory_arlen + 1;
  wire [41-1:0] pack_read_req_packed_20;
  assign pack_read_req_packed_20 = { pack_read_req_global_addr_18, pack_read_req_size_19 };
  assign _memory_rreq_fifo_wdata = ((_memory_raddr_fsm == 1) && memory_arvalid && memory_arready)? pack_read_req_packed_20 : 'hx;
  assign _memory_rreq_fifo_enq = ((_memory_raddr_fsm == 1) && memory_arvalid && memory_arready)? (_memory_raddr_fsm == 1) && memory_arvalid && memory_arready && !_memory_rreq_fifo_almost_full : 0;
  localparam _tmp_21 = 1;
  wire [_tmp_21-1:0] _tmp_22;
  assign _tmp_22 = !_memory_rreq_fifo_almost_full;
  reg [_tmp_21-1:0] __tmp_22_1;
  wire [32-1:0] unpack_read_req_global_addr_23;
  wire [9-1:0] unpack_read_req_size_24;
  assign unpack_read_req_global_addr_23 = _memory_rreq_fifo_rdata[40:9];
  assign unpack_read_req_size_24 = _memory_rreq_fifo_rdata[8:0];
  assign _memory_rreq_fifo_deq = ((_memory_rdata_fsm == 0) && !_memory_rreq_fifo_empty && !_memory_rreq_fifo_empty)? 1 : 0;
  reg [32-1:0] _d1__memory_rdata_fsm;
  reg __memory_rdata_fsm_cond_11_0_1;
  assign memory_awaddr = maxi_awaddr;
  assign memory_awlen = maxi_awlen;
  assign memory_awsize = maxi_awsize;
  assign memory_awburst = maxi_awburst;
  assign memory_awlock = maxi_awlock;
  assign memory_awcache = maxi_awcache;
  assign memory_awprot = maxi_awprot;
  assign memory_awqos = maxi_awqos;
  assign memory_awuser = maxi_awuser;
  assign memory_awvalid = maxi_awvalid;
  wire _tmp_25;
  assign _tmp_25 = memory_awready;

  always @(*) begin
    maxi_awready = _tmp_25;
  end

  assign memory_wdata = maxi_wdata;
  assign memory_wstrb = maxi_wstrb;
  assign memory_wlast = maxi_wlast;
  assign memory_wvalid = maxi_wvalid;
  wire _tmp_26;
  assign _tmp_26 = memory_wready;

  always @(*) begin
    maxi_wready = _tmp_26;
  end

  wire [2-1:0] _tmp_27;
  assign _tmp_27 = memory_bresp;

  always @(*) begin
    maxi_bresp = _tmp_27;
  end

  wire _tmp_28;
  assign _tmp_28 = memory_bvalid;

  always @(*) begin
    maxi_bvalid = _tmp_28;
  end

  assign memory_bready = maxi_bready;
  assign memory_araddr = maxi_araddr;
  assign memory_arlen = maxi_arlen;
  assign memory_arsize = maxi_arsize;
  assign memory_arburst = maxi_arburst;
  assign memory_arlock = maxi_arlock;
  assign memory_arcache = maxi_arcache;
  assign memory_arprot = maxi_arprot;
  assign memory_arqos = maxi_arqos;
  assign memory_aruser = maxi_aruser;
  assign memory_arvalid = maxi_arvalid;
  wire _tmp_29;
  assign _tmp_29 = memory_arready;

  always @(*) begin
    maxi_arready = _tmp_29;
  end

  wire [32-1:0] _tmp_30;
  assign _tmp_30 = memory_rdata;

  always @(*) begin
    maxi_rdata = _tmp_30;
  end

  wire [2-1:0] _tmp_31;
  assign _tmp_31 = memory_rresp;

  always @(*) begin
    maxi_rresp = _tmp_31;
  end

  wire _tmp_32;
  assign _tmp_32 = memory_rlast;

  always @(*) begin
    maxi_rlast = _tmp_32;
  end

  wire _tmp_33;
  assign _tmp_33 = memory_rvalid;

  always @(*) begin
    maxi_rvalid = _tmp_33;
  end

  assign memory_rready = maxi_rready;
  reg [32-1:0] _saxi_awaddr;
  wire [4-1:0] _saxi_awcache;
  wire [3-1:0] _saxi_awprot;
  reg _saxi_awvalid;
  wire _saxi_awready;
  assign _saxi_awcache = 3;
  assign _saxi_awprot = 0;
  wire [32-1:0] _saxi_wdata;
  wire [4-1:0] _saxi_wstrb;
  wire _saxi_wvalid;
  wire _saxi_wready;
  reg [32-1:0] __saxi_wdata_sb_0;
  reg [4-1:0] __saxi_wstrb_sb_0;
  reg __saxi_wvalid_sb_0;
  wire __saxi_wready_sb_0;
  wire [4-1:0] _sb__saxi_writedata_s_value_34;
  assign _sb__saxi_writedata_s_value_34 = __saxi_wstrb_sb_0;
  wire [32-1:0] _sb__saxi_writedata_s_value_35;
  assign _sb__saxi_writedata_s_value_35 = __saxi_wdata_sb_0;
  wire [36-1:0] _sb__saxi_writedata_s_data_36;
  assign _sb__saxi_writedata_s_data_36 = { _sb__saxi_writedata_s_value_34, _sb__saxi_writedata_s_value_35 };
  wire _sb__saxi_writedata_s_valid_37;
  assign _sb__saxi_writedata_s_valid_37 = __saxi_wvalid_sb_0;
  wire _sb__saxi_writedata_m_ready_38;
  assign _sb__saxi_writedata_m_ready_38 = _saxi_wready;
  reg [36-1:0] _sb__saxi_writedata_data_39;
  reg _sb__saxi_writedata_valid_40;
  wire _sb__saxi_writedata_ready_41;
  reg [36-1:0] _sb__saxi_writedata_tmp_data_42;
  reg _sb__saxi_writedata_tmp_valid_43;
  wire [36-1:0] _sb__saxi_writedata_next_data_44;
  wire _sb__saxi_writedata_next_valid_45;
  assign _sb__saxi_writedata_ready_41 = !_sb__saxi_writedata_tmp_valid_43;
  assign _sb__saxi_writedata_next_data_44 = (_sb__saxi_writedata_tmp_valid_43)? _sb__saxi_writedata_tmp_data_42 : _sb__saxi_writedata_s_data_36;
  assign _sb__saxi_writedata_next_valid_45 = _sb__saxi_writedata_tmp_valid_43 || _sb__saxi_writedata_s_valid_37;
  wire [4-1:0] _sb__saxi_writedata_m_value_46;
  assign _sb__saxi_writedata_m_value_46 = _sb__saxi_writedata_data_39[35:32];
  wire [32-1:0] _sb__saxi_writedata_m_value_47;
  assign _sb__saxi_writedata_m_value_47 = _sb__saxi_writedata_data_39[31:0];
  assign __saxi_wready_sb_0 = _sb__saxi_writedata_ready_41;
  assign _saxi_wdata = _sb__saxi_writedata_m_value_47;
  assign _saxi_wstrb = _sb__saxi_writedata_m_value_46;
  assign _saxi_wvalid = _sb__saxi_writedata_valid_40;
  wire [2-1:0] _saxi_bresp;
  wire _saxi_bvalid;
  wire _saxi_bready;
  assign _saxi_bready = 1;
  reg [32-1:0] _saxi_araddr;
  wire [4-1:0] _saxi_arcache;
  wire [3-1:0] _saxi_arprot;
  reg _saxi_arvalid;
  wire _saxi_arready;
  assign _saxi_arcache = 3;
  assign _saxi_arprot = 0;
  wire [32-1:0] _saxi_rdata;
  wire [2-1:0] _saxi_rresp;
  wire _saxi_rvalid;
  wire _saxi_rready;
  wire [32-1:0] __saxi_rdata_sb_0;
  wire __saxi_rvalid_sb_0;
  wire __saxi_rready_sb_0;
  wire [32-1:0] _sb__saxi_readdata_s_value_48;
  assign _sb__saxi_readdata_s_value_48 = _saxi_rdata;
  wire [32-1:0] _sb__saxi_readdata_s_data_49;
  assign _sb__saxi_readdata_s_data_49 = { _sb__saxi_readdata_s_value_48 };
  wire _sb__saxi_readdata_s_valid_50;
  assign _sb__saxi_readdata_s_valid_50 = _saxi_rvalid;
  wire _sb__saxi_readdata_m_ready_51;
  assign _sb__saxi_readdata_m_ready_51 = __saxi_rready_sb_0;
  reg [32-1:0] _sb__saxi_readdata_data_52;
  reg _sb__saxi_readdata_valid_53;
  wire _sb__saxi_readdata_ready_54;
  reg [32-1:0] _sb__saxi_readdata_tmp_data_55;
  reg _sb__saxi_readdata_tmp_valid_56;
  wire [32-1:0] _sb__saxi_readdata_next_data_57;
  wire _sb__saxi_readdata_next_valid_58;
  assign _sb__saxi_readdata_ready_54 = !_sb__saxi_readdata_tmp_valid_56;
  assign _sb__saxi_readdata_next_data_57 = (_sb__saxi_readdata_tmp_valid_56)? _sb__saxi_readdata_tmp_data_55 : _sb__saxi_readdata_s_data_49;
  assign _sb__saxi_readdata_next_valid_58 = _sb__saxi_readdata_tmp_valid_56 || _sb__saxi_readdata_s_valid_50;
  wire [32-1:0] _sb__saxi_readdata_m_value_59;
  assign _sb__saxi_readdata_m_value_59 = _sb__saxi_readdata_data_52[31:0];
  assign __saxi_rdata_sb_0 = _sb__saxi_readdata_m_value_59;
  assign __saxi_rvalid_sb_0 = _sb__saxi_readdata_valid_53;
  assign _saxi_rready = _sb__saxi_readdata_ready_54;
  reg [3-1:0] __saxi_outstanding_wcount;
  wire __saxi_has_outstanding_write;
  assign __saxi_has_outstanding_write = (__saxi_outstanding_wcount > 0) || _saxi_awvalid;
  wire [32-1:0] _tmp_60;
  assign _tmp_60 = _saxi_awaddr;

  always @(*) begin
    saxi_awaddr = _tmp_60;
  end

  wire [4-1:0] _tmp_61;
  assign _tmp_61 = _saxi_awcache;

  always @(*) begin
    saxi_awcache = _tmp_61;
  end

  wire [3-1:0] _tmp_62;
  assign _tmp_62 = _saxi_awprot;

  always @(*) begin
    saxi_awprot = _tmp_62;
  end

  wire _tmp_63;
  assign _tmp_63 = _saxi_awvalid;

  always @(*) begin
    saxi_awvalid = _tmp_63;
  end

  assign _saxi_awready = saxi_awready;
  wire [32-1:0] _tmp_64;
  assign _tmp_64 = _saxi_wdata;

  always @(*) begin
    saxi_wdata = _tmp_64;
  end

  wire [4-1:0] _tmp_65;
  assign _tmp_65 = _saxi_wstrb;

  always @(*) begin
    saxi_wstrb = _tmp_65;
  end

  wire _tmp_66;
  assign _tmp_66 = _saxi_wvalid;

  always @(*) begin
    saxi_wvalid = _tmp_66;
  end

  assign _saxi_wready = saxi_wready;
  assign _saxi_bresp = saxi_bresp;
  assign _saxi_bvalid = saxi_bvalid;
  wire _tmp_67;
  assign _tmp_67 = _saxi_bready;

  always @(*) begin
    saxi_bready = _tmp_67;
  end

  wire [32-1:0] _tmp_68;
  assign _tmp_68 = _saxi_araddr;

  always @(*) begin
    saxi_araddr = _tmp_68;
  end

  wire [4-1:0] _tmp_69;
  assign _tmp_69 = _saxi_arcache;

  always @(*) begin
    saxi_arcache = _tmp_69;
  end

  wire [3-1:0] _tmp_70;
  assign _tmp_70 = _saxi_arprot;

  always @(*) begin
    saxi_arprot = _tmp_70;
  end

  wire _tmp_71;
  assign _tmp_71 = _saxi_arvalid;

  always @(*) begin
    saxi_arvalid = _tmp_71;
  end

  assign _saxi_arready = saxi_arready;
  assign _saxi_rdata = saxi_rdata;
  assign _saxi_rresp = saxi_rresp;
  assign _saxi_rvalid = saxi_rvalid;
  wire _tmp_72;
  assign _tmp_72 = _saxi_rready;

  always @(*) begin
    saxi_rready = _tmp_72;
  end

  reg [32-1:0] time_counter;
  reg [32-1:0] th_ctrl;
  localparam th_ctrl_init = 0;
  reg signed [32-1:0] _th_ctrl_i_0;
  reg __saxi_waddr_cond_0_1;
  reg __saxi_wdata_cond_0_1;
  reg signed [32-1:0] _th_ctrl_start_time_1;
  reg __saxi_waddr_cond_1_1;
  reg __saxi_wdata_cond_1_1;
  reg __saxi_raddr_cond_0_1;
  reg signed [32-1:0] axim_rdata_73;
  reg __saxi_raddr_cond_1_1;
  reg signed [32-1:0] axim_rdata_74;
  assign __saxi_rready_sb_0 = (th_ctrl == 17) || (th_ctrl == 22);
  reg signed [32-1:0] _th_ctrl_end_time_2;
  reg signed [32-1:0] _th_ctrl_ok_3;
  reg signed [32-1:0] _th_ctrl_bat_4;
  reg signed [32-1:0] _th_ctrl_x_5;
  reg signed [16-1:0] rdata_75;
  reg signed [32-1:0] _th_ctrl_orig_6;
  reg signed [16-1:0] rdata_76;
  reg signed [32-1:0] _th_ctrl_check_7;

  hello_nngen
  uut
  (
    .CLK(CLK),
    .RESETN(RESETN),
    .irq(irq),
    .maxi_awaddr(maxi_awaddr),
    .maxi_awlen(maxi_awlen),
    .maxi_awsize(maxi_awsize),
    .maxi_awburst(maxi_awburst),
    .maxi_awlock(maxi_awlock),
    .maxi_awcache(maxi_awcache),
    .maxi_awprot(maxi_awprot),
    .maxi_awqos(maxi_awqos),
    .maxi_awuser(maxi_awuser),
    .maxi_awvalid(maxi_awvalid),
    .maxi_awready(maxi_awready),
    .maxi_wdata(maxi_wdata),
    .maxi_wstrb(maxi_wstrb),
    .maxi_wlast(maxi_wlast),
    .maxi_wvalid(maxi_wvalid),
    .maxi_wready(maxi_wready),
    .maxi_bresp(maxi_bresp),
    .maxi_bvalid(maxi_bvalid),
    .maxi_bready(maxi_bready),
    .maxi_araddr(maxi_araddr),
    .maxi_arlen(maxi_arlen),
    .maxi_arsize(maxi_arsize),
    .maxi_arburst(maxi_arburst),
    .maxi_arlock(maxi_arlock),
    .maxi_arcache(maxi_arcache),
    .maxi_arprot(maxi_arprot),
    .maxi_arqos(maxi_arqos),
    .maxi_aruser(maxi_aruser),
    .maxi_arvalid(maxi_arvalid),
    .maxi_arready(maxi_arready),
    .maxi_rdata(maxi_rdata),
    .maxi_rresp(maxi_rresp),
    .maxi_rlast(maxi_rlast),
    .maxi_rvalid(maxi_rvalid),
    .maxi_rready(maxi_rready),
    .saxi_awaddr(saxi_awaddr),
    .saxi_awcache(saxi_awcache),
    .saxi_awprot(saxi_awprot),
    .saxi_awvalid(saxi_awvalid),
    .saxi_awready(saxi_awready),
    .saxi_wdata(saxi_wdata),
    .saxi_wstrb(saxi_wstrb),
    .saxi_wvalid(saxi_wvalid),
    .saxi_wready(saxi_wready),
    .saxi_bresp(saxi_bresp),
    .saxi_bvalid(saxi_bvalid),
    .saxi_bready(saxi_bready),
    .saxi_araddr(saxi_araddr),
    .saxi_arcache(saxi_arcache),
    .saxi_arprot(saxi_arprot),
    .saxi_arvalid(saxi_arvalid),
    .saxi_arready(saxi_arready),
    .saxi_rdata(saxi_rdata),
    .saxi_rresp(saxi_rresp),
    .saxi_rvalid(saxi_rvalid),
    .saxi_rready(saxi_rready)
  );


  initial begin
    CLK = 0;
    forever begin
      #5 CLK = !CLK;
    end
  end


  initial begin
    RESETN = 1;
    memory_awready = 0;
    memory_bvalid = 0;
    memory_arready = 0;
    memory_rdata = 0;
    memory_rlast = 0;
    memory_rvalid = 0;
    _memory_waddr_fsm = _memory_waddr_fsm_init;
    _memory_wdata_fsm = _memory_wdata_fsm_init;
    _memory_raddr_fsm = _memory_raddr_fsm_init;
    _memory_rdata_fsm = _memory_rdata_fsm_init;
    count__memory_wreq_fifo = 0;
    count__memory_rreq_fifo = 0;
    count__memory_wdata_fifo = 0;
    __tmp_5_1 = 0;
    _write_count = 0;
    _write_addr = 0;
    _read_count = 0;
    _read_addr = 0;
    _sleep_interval_count = 0;
    _keep_sleep_count = 0;
    __tmp_10_1 = 0;
    __tmp_22_1 = 0;
    _d1__memory_rdata_fsm = _memory_rdata_fsm_init;
    __memory_rdata_fsm_cond_11_0_1 = 0;
    _saxi_awaddr = 0;
    _saxi_awvalid = 0;
    __saxi_wdata_sb_0 = 0;
    __saxi_wstrb_sb_0 = 0;
    __saxi_wvalid_sb_0 = 0;
    _sb__saxi_writedata_data_39 = 0;
    _sb__saxi_writedata_valid_40 = 0;
    _sb__saxi_writedata_tmp_data_42 = 0;
    _sb__saxi_writedata_tmp_valid_43 = 0;
    _saxi_araddr = 0;
    _saxi_arvalid = 0;
    _sb__saxi_readdata_data_52 = 0;
    _sb__saxi_readdata_valid_53 = 0;
    _sb__saxi_readdata_tmp_data_55 = 0;
    _sb__saxi_readdata_tmp_valid_56 = 0;
    __saxi_outstanding_wcount = 0;
    time_counter = 0;
    th_ctrl = th_ctrl_init;
    _th_ctrl_i_0 = 0;
    __saxi_waddr_cond_0_1 = 0;
    __saxi_wdata_cond_0_1 = 0;
    _th_ctrl_start_time_1 = 0;
    __saxi_waddr_cond_1_1 = 0;
    __saxi_wdata_cond_1_1 = 0;
    __saxi_raddr_cond_0_1 = 0;
    axim_rdata_73 = 0;
    __saxi_raddr_cond_1_1 = 0;
    axim_rdata_74 = 0;
    _th_ctrl_end_time_2 = 0;
    _th_ctrl_ok_3 = 0;
    _th_ctrl_bat_4 = 0;
    _th_ctrl_x_5 = 0;
    rdata_75 = 0;
    _th_ctrl_orig_6 = 0;
    rdata_76 = 0;
    _th_ctrl_check_7 = 0;
    #100;
    RESETN = 0;
    #100;
    RESETN = 1;
    #10000000;
    $finish;
  end


  always @(posedge CLK) begin
    if(RST) begin
      _keep_sleep_count <= 0;
      _sleep_interval_count <= 0;
    end else begin
      if(_sleep_interval_count == 15) begin
        _keep_sleep_count <= _keep_sleep_count + 1;
      end 
      if((_sleep_interval_count == 15) && (_keep_sleep_count == 3)) begin
        _keep_sleep_count <= 0;
      end 
      if(_sleep_interval_count < 15) begin
        _sleep_interval_count <= _sleep_interval_count + 1;
      end 
      if((_keep_sleep_count == 3) && (_sleep_interval_count == 15)) begin
        _sleep_interval_count <= 0;
      end 
      if((_memory_wdata_fsm == 1) && write_data_wvalid_16 && write_data_wready_17 && pack_write_data_wstrb_14[0]) begin
        _memory_mem[_write_addr + 0] <= pack_write_data_wdata_13[7:0];
      end 
      if((_memory_wdata_fsm == 1) && write_data_wvalid_16 && write_data_wready_17 && pack_write_data_wstrb_14[1]) begin
        _memory_mem[_write_addr + 1] <= pack_write_data_wdata_13[15:8];
      end 
      if((_memory_wdata_fsm == 1) && write_data_wvalid_16 && write_data_wready_17 && pack_write_data_wstrb_14[2]) begin
        _memory_mem[_write_addr + 2] <= pack_write_data_wdata_13[23:16];
      end 
      if((_memory_wdata_fsm == 1) && write_data_wvalid_16 && write_data_wready_17 && pack_write_data_wstrb_14[3]) begin
        _memory_mem[_write_addr + 3] <= pack_write_data_wdata_13[31:24];
      end 
    end
  end

  localparam _memory_waddr_fsm_1 = 1;
  localparam _memory_waddr_fsm_2 = 2;
  localparam _memory_waddr_fsm_3 = 3;
  localparam _memory_waddr_fsm_4 = 4;
  localparam _memory_waddr_fsm_5 = 5;
  localparam _memory_waddr_fsm_6 = 6;
  localparam _memory_waddr_fsm_7 = 7;
  localparam _memory_waddr_fsm_8 = 8;
  localparam _memory_waddr_fsm_9 = 9;
  localparam _memory_waddr_fsm_10 = 10;
  localparam _memory_waddr_fsm_11 = 11;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_waddr_fsm <= _memory_waddr_fsm_init;
      memory_awready <= 0;
    end else begin
      case(_memory_waddr_fsm)
        _memory_waddr_fsm_init: begin
          memory_awready <= 0;
          if(memory_awvalid) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_1;
          end 
        end
        _memory_waddr_fsm_1: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_2;
        end
        _memory_waddr_fsm_2: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_3;
        end
        _memory_waddr_fsm_3: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_4;
        end
        _memory_waddr_fsm_4: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_5;
        end
        _memory_waddr_fsm_5: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_6;
        end
        _memory_waddr_fsm_6: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_7;
        end
        _memory_waddr_fsm_7: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_8;
        end
        _memory_waddr_fsm_8: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_9;
        end
        _memory_waddr_fsm_9: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_10;
        end
        _memory_waddr_fsm_10: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_11;
        end
        _memory_waddr_fsm_11: begin
          if(!_memory_wreq_fifo_almost_full) begin
            memory_awready <= 1;
          end 
          if(memory_awvalid && memory_awready) begin
            memory_awready <= 0;
          end 
          if(!memory_awvalid) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_init;
          end 
          if(memory_awvalid && memory_awready) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_wdata_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_wdata_fsm <= _memory_wdata_fsm_init;
      memory_bvalid <= 0;
      _write_addr <= 0;
      _write_count <= 0;
    end else begin
      case(_memory_wdata_fsm)
        _memory_wdata_fsm_init: begin
          memory_bvalid <= 0;
          if(!_memory_wreq_fifo_empty) begin
            _write_addr <= unpack_write_req_global_addr_11;
            _write_count <= unpack_write_req_size_12;
          end 
          if(!_memory_wreq_fifo_empty) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_1;
          end 
        end
        _memory_wdata_fsm_1: begin
          if(write_data_wvalid_16 && write_data_wready_17) begin
            _write_addr <= _write_addr + 4;
            _write_count <= _write_count - 1;
          end 
          if(write_data_wvalid_16 && write_data_wready_17 && (_write_count == 1)) begin
            memory_bvalid <= 1;
          end 
          if(write_data_wvalid_16 && write_data_wready_17 && pack_write_data_wlast_15) begin
            memory_bvalid <= 1;
          end 
          if(write_data_wvalid_16 && write_data_wready_17 && (_write_count == 1)) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_init;
          end 
          if(write_data_wvalid_16 && write_data_wready_17 && pack_write_data_wlast_15) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_raddr_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_raddr_fsm <= _memory_raddr_fsm_init;
      memory_arready <= 0;
    end else begin
      case(_memory_raddr_fsm)
        _memory_raddr_fsm_init: begin
          memory_arready <= 0;
          if(memory_arvalid) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_1;
          end 
        end
        _memory_raddr_fsm_1: begin
          if(!_memory_rreq_fifo_almost_full) begin
            memory_arready <= 1;
          end 
          if(memory_arvalid && memory_arready) begin
            memory_arready <= 0;
          end 
          if(!memory_arvalid) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_init;
          end 
          if(memory_arvalid && memory_arready) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_rdata_fsm_1 = 1;
  localparam _memory_rdata_fsm_2 = 2;
  localparam _memory_rdata_fsm_3 = 3;
  localparam _memory_rdata_fsm_4 = 4;
  localparam _memory_rdata_fsm_5 = 5;
  localparam _memory_rdata_fsm_6 = 6;
  localparam _memory_rdata_fsm_7 = 7;
  localparam _memory_rdata_fsm_8 = 8;
  localparam _memory_rdata_fsm_9 = 9;
  localparam _memory_rdata_fsm_10 = 10;
  localparam _memory_rdata_fsm_11 = 11;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_rdata_fsm <= _memory_rdata_fsm_init;
      _d1__memory_rdata_fsm <= _memory_rdata_fsm_init;
      _read_addr <= 0;
      _read_count <= 0;
      memory_rdata[7:0] <= (0 >> 0) & { 8{ 1'd1 } };
      memory_rdata[15:8] <= (0 >> 8) & { 8{ 1'd1 } };
      memory_rdata[23:16] <= (0 >> 16) & { 8{ 1'd1 } };
      memory_rdata[31:24] <= (0 >> 24) & { 8{ 1'd1 } };
      memory_rvalid <= 0;
      memory_rlast <= 0;
      __memory_rdata_fsm_cond_11_0_1 <= 0;
      memory_rdata <= 0;
    end else begin
      _d1__memory_rdata_fsm <= _memory_rdata_fsm;
      case(_d1__memory_rdata_fsm)
        _memory_rdata_fsm_11: begin
          if(__memory_rdata_fsm_cond_11_0_1) begin
            memory_rvalid <= 0;
            memory_rlast <= 0;
          end 
        end
      endcase
      case(_memory_rdata_fsm)
        _memory_rdata_fsm_init: begin
          if(!_memory_rreq_fifo_empty) begin
            _read_addr <= unpack_read_req_global_addr_23;
            _read_count <= unpack_read_req_size_24;
          end 
          if(!_memory_rreq_fifo_empty) begin
            _memory_rdata_fsm <= _memory_rdata_fsm_1;
          end 
        end
        _memory_rdata_fsm_1: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_2;
        end
        _memory_rdata_fsm_2: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_3;
        end
        _memory_rdata_fsm_3: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_4;
        end
        _memory_rdata_fsm_4: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_5;
        end
        _memory_rdata_fsm_5: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_6;
        end
        _memory_rdata_fsm_6: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_7;
        end
        _memory_rdata_fsm_7: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_8;
        end
        _memory_rdata_fsm_8: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_9;
        end
        _memory_rdata_fsm_9: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_10;
        end
        _memory_rdata_fsm_10: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_11;
        end
        _memory_rdata_fsm_11: begin
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[7:0] <= _memory_mem[_read_addr + 0];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[15:8] <= _memory_mem[_read_addr + 1];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[23:16] <= _memory_mem[_read_addr + 2];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[31:24] <= _memory_mem[_read_addr + 3];
          end 
          if((_sleep_interval_count < 15) && (_read_count > 0) && memory_rready | !memory_rvalid) begin
            memory_rvalid <= 1;
            _read_addr <= _read_addr + 4;
            _read_count <= _read_count - 1;
          end 
          if((_sleep_interval_count < 15) && (_read_count == 1) && memory_rready | !memory_rvalid) begin
            memory_rlast <= 1;
          end 
          __memory_rdata_fsm_cond_11_0_1 <= 1;
          if(memory_rvalid && !memory_rready) begin
            memory_rvalid <= memory_rvalid;
            memory_rdata <= memory_rdata;
            memory_rlast <= memory_rlast;
          end 
          if(memory_rvalid && memory_rready && (_read_count == 0)) begin
            _memory_rdata_fsm <= _memory_rdata_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__memory_wreq_fifo <= 0;
      __tmp_10_1 <= 0;
    end else begin
      if(_memory_wreq_fifo_enq && !_memory_wreq_fifo_full && (_memory_wreq_fifo_deq && !_memory_wreq_fifo_empty)) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo;
      end else if(_memory_wreq_fifo_enq && !_memory_wreq_fifo_full) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo + 1;
      end else if(_memory_wreq_fifo_deq && !_memory_wreq_fifo_empty) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo - 1;
      end 
      __tmp_10_1 <= _tmp_10;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__memory_rreq_fifo <= 0;
      __tmp_22_1 <= 0;
    end else begin
      if(_memory_rreq_fifo_enq && !_memory_rreq_fifo_full && (_memory_rreq_fifo_deq && !_memory_rreq_fifo_empty)) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo;
      end else if(_memory_rreq_fifo_enq && !_memory_rreq_fifo_full) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo + 1;
      end else if(_memory_rreq_fifo_deq && !_memory_rreq_fifo_empty) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo - 1;
      end 
      __tmp_22_1 <= _tmp_22;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__memory_wdata_fifo <= 0;
      __tmp_5_1 <= 0;
    end else begin
      if(_memory_wdata_fifo_enq && !_memory_wdata_fifo_full && (_memory_wdata_fifo_deq && !_memory_wdata_fifo_empty)) begin
        count__memory_wdata_fifo <= count__memory_wdata_fifo;
      end else if(_memory_wdata_fifo_enq && !_memory_wdata_fifo_full) begin
        count__memory_wdata_fifo <= count__memory_wdata_fifo + 1;
      end else if(_memory_wdata_fifo_deq && !_memory_wdata_fifo_empty) begin
        count__memory_wdata_fifo <= count__memory_wdata_fifo - 1;
      end 
      __tmp_5_1 <= _tmp_5;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _saxi_awaddr <= 0;
      _saxi_awvalid <= 0;
      __saxi_waddr_cond_0_1 <= 0;
      __saxi_waddr_cond_1_1 <= 0;
    end else begin
      if(__saxi_waddr_cond_0_1) begin
        _saxi_awvalid <= 0;
      end 
      if(__saxi_waddr_cond_1_1) begin
        _saxi_awvalid <= 0;
      end 
      if((th_ctrl == 4) && ((__saxi_outstanding_wcount == 0) && (_saxi_awready || !_saxi_awvalid))) begin
        _saxi_awaddr <= 132;
        _saxi_awvalid <= 1;
      end 
      __saxi_waddr_cond_0_1 <= 1;
      if(_saxi_awvalid && !_saxi_awready) begin
        _saxi_awvalid <= _saxi_awvalid;
      end 
      if((th_ctrl == 10) && ((__saxi_outstanding_wcount == 0) && (_saxi_awready || !_saxi_awvalid))) begin
        _saxi_awaddr <= 16;
        _saxi_awvalid <= 1;
      end 
      __saxi_waddr_cond_1_1 <= 1;
      if(_saxi_awvalid && !_saxi_awready) begin
        _saxi_awvalid <= _saxi_awvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __saxi_wdata_sb_0 <= 0;
      __saxi_wvalid_sb_0 <= 0;
      __saxi_wstrb_sb_0 <= 0;
      __saxi_wdata_cond_0_1 <= 0;
      __saxi_wdata_cond_1_1 <= 0;
    end else begin
      if(__saxi_wdata_cond_0_1) begin
        __saxi_wvalid_sb_0 <= 0;
      end 
      if(__saxi_wdata_cond_1_1) begin
        __saxi_wvalid_sb_0 <= 0;
      end 
      if((th_ctrl == 6) && (__saxi_wready_sb_0 || !__saxi_wvalid_sb_0)) begin
        __saxi_wdata_sb_0 <= 8482048;
        __saxi_wvalid_sb_0 <= 1;
        __saxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      __saxi_wdata_cond_0_1 <= 1;
      if(__saxi_wvalid_sb_0 && !__saxi_wready_sb_0) begin
        __saxi_wvalid_sb_0 <= __saxi_wvalid_sb_0;
      end 
      if((th_ctrl == 12) && (__saxi_wready_sb_0 || !__saxi_wvalid_sb_0)) begin
        __saxi_wdata_sb_0 <= 1;
        __saxi_wvalid_sb_0 <= 1;
        __saxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      __saxi_wdata_cond_1_1 <= 1;
      if(__saxi_wvalid_sb_0 && !__saxi_wready_sb_0) begin
        __saxi_wvalid_sb_0 <= __saxi_wvalid_sb_0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _sb__saxi_writedata_data_39 <= 0;
      _sb__saxi_writedata_valid_40 <= 0;
      _sb__saxi_writedata_tmp_data_42 <= 0;
      _sb__saxi_writedata_tmp_valid_43 <= 0;
    end else begin
      if(_sb__saxi_writedata_m_ready_38 || !_sb__saxi_writedata_valid_40) begin
        _sb__saxi_writedata_data_39 <= _sb__saxi_writedata_next_data_44;
        _sb__saxi_writedata_valid_40 <= _sb__saxi_writedata_next_valid_45;
      end 
      if(!_sb__saxi_writedata_tmp_valid_43 && _sb__saxi_writedata_valid_40 && !_sb__saxi_writedata_m_ready_38) begin
        _sb__saxi_writedata_tmp_data_42 <= _sb__saxi_writedata_s_data_36;
        _sb__saxi_writedata_tmp_valid_43 <= _sb__saxi_writedata_s_valid_37;
      end 
      if(_sb__saxi_writedata_tmp_valid_43 && _sb__saxi_writedata_m_ready_38) begin
        _sb__saxi_writedata_tmp_valid_43 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _saxi_araddr <= 0;
      _saxi_arvalid <= 0;
      __saxi_raddr_cond_0_1 <= 0;
      __saxi_raddr_cond_1_1 <= 0;
    end else begin
      if(__saxi_raddr_cond_0_1) begin
        _saxi_arvalid <= 0;
      end 
      if(__saxi_raddr_cond_1_1) begin
        _saxi_arvalid <= 0;
      end 
      if((th_ctrl == 15) && (_saxi_arready || !_saxi_arvalid)) begin
        _saxi_araddr <= 16;
        _saxi_arvalid <= 1;
      end 
      __saxi_raddr_cond_0_1 <= 1;
      if(_saxi_arvalid && !_saxi_arready) begin
        _saxi_arvalid <= _saxi_arvalid;
      end 
      if((th_ctrl == 20) && (_saxi_arready || !_saxi_arvalid)) begin
        _saxi_araddr <= 20;
        _saxi_arvalid <= 1;
      end 
      __saxi_raddr_cond_1_1 <= 1;
      if(_saxi_arvalid && !_saxi_arready) begin
        _saxi_arvalid <= _saxi_arvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _sb__saxi_readdata_data_52 <= 0;
      _sb__saxi_readdata_valid_53 <= 0;
      _sb__saxi_readdata_tmp_data_55 <= 0;
      _sb__saxi_readdata_tmp_valid_56 <= 0;
    end else begin
      if(_sb__saxi_readdata_m_ready_51 || !_sb__saxi_readdata_valid_53) begin
        _sb__saxi_readdata_data_52 <= _sb__saxi_readdata_next_data_57;
        _sb__saxi_readdata_valid_53 <= _sb__saxi_readdata_next_valid_58;
      end 
      if(!_sb__saxi_readdata_tmp_valid_56 && _sb__saxi_readdata_valid_53 && !_sb__saxi_readdata_m_ready_51) begin
        _sb__saxi_readdata_tmp_data_55 <= _sb__saxi_readdata_s_data_49;
        _sb__saxi_readdata_tmp_valid_56 <= _sb__saxi_readdata_s_valid_50;
      end 
      if(_sb__saxi_readdata_tmp_valid_56 && _sb__saxi_readdata_m_ready_51) begin
        _sb__saxi_readdata_tmp_valid_56 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __saxi_outstanding_wcount <= 0;
    end else begin
      if(_saxi_awvalid && _saxi_awready && !(_saxi_bvalid && _saxi_bready) && (__saxi_outstanding_wcount < 7)) begin
        __saxi_outstanding_wcount <= __saxi_outstanding_wcount + 1;
      end 
      if(!(_saxi_awvalid && _saxi_awready) && (_saxi_bvalid && _saxi_bready) && (__saxi_outstanding_wcount > 0)) begin
        __saxi_outstanding_wcount <= __saxi_outstanding_wcount - 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      time_counter <= 0;
    end else begin
      time_counter <= time_counter + 1;
    end
  end

  localparam th_ctrl_1 = 1;
  localparam th_ctrl_2 = 2;
  localparam th_ctrl_3 = 3;
  localparam th_ctrl_4 = 4;
  localparam th_ctrl_5 = 5;
  localparam th_ctrl_6 = 6;
  localparam th_ctrl_7 = 7;
  localparam th_ctrl_8 = 8;
  localparam th_ctrl_9 = 9;
  localparam th_ctrl_10 = 10;
  localparam th_ctrl_11 = 11;
  localparam th_ctrl_12 = 12;
  localparam th_ctrl_13 = 13;
  localparam th_ctrl_14 = 14;
  localparam th_ctrl_15 = 15;
  localparam th_ctrl_16 = 16;
  localparam th_ctrl_17 = 17;
  localparam th_ctrl_18 = 18;
  localparam th_ctrl_19 = 19;
  localparam th_ctrl_20 = 20;
  localparam th_ctrl_21 = 21;
  localparam th_ctrl_22 = 22;
  localparam th_ctrl_23 = 23;
  localparam th_ctrl_24 = 24;
  localparam th_ctrl_25 = 25;
  localparam th_ctrl_26 = 26;
  localparam th_ctrl_27 = 27;
  localparam th_ctrl_28 = 28;
  localparam th_ctrl_29 = 29;
  localparam th_ctrl_30 = 30;
  localparam th_ctrl_31 = 31;
  localparam th_ctrl_32 = 32;
  localparam th_ctrl_33 = 33;
  localparam th_ctrl_34 = 34;
  localparam th_ctrl_35 = 35;
  localparam th_ctrl_36 = 36;
  localparam th_ctrl_37 = 37;
  localparam th_ctrl_38 = 38;
  localparam th_ctrl_39 = 39;
  localparam th_ctrl_40 = 40;
  localparam th_ctrl_41 = 41;
  localparam th_ctrl_42 = 42;
  localparam th_ctrl_43 = 43;
  localparam th_ctrl_44 = 44;
  localparam th_ctrl_45 = 45;
  localparam th_ctrl_46 = 46;
  localparam th_ctrl_47 = 47;
  localparam th_ctrl_48 = 48;

  always @(posedge CLK) begin
    if(RST) begin
      th_ctrl <= th_ctrl_init;
      _th_ctrl_i_0 <= 0;
      _th_ctrl_start_time_1 <= 0;
      axim_rdata_73 <= 0;
      axim_rdata_74 <= 0;
      _th_ctrl_end_time_2 <= 0;
      _th_ctrl_ok_3 <= 0;
      _th_ctrl_bat_4 <= 0;
      _th_ctrl_x_5 <= 0;
      rdata_75 <= 0;
      _th_ctrl_orig_6 <= 0;
      rdata_76 <= 0;
      _th_ctrl_check_7 <= 0;
    end else begin
      case(th_ctrl)
        th_ctrl_init: begin
          th_ctrl <= th_ctrl_1;
        end
        th_ctrl_1: begin
          _th_ctrl_i_0 <= 0;
          th_ctrl <= th_ctrl_2;
        end
        th_ctrl_2: begin
          if(_th_ctrl_i_0 < 100) begin
            th_ctrl <= th_ctrl_3;
          end else begin
            th_ctrl <= th_ctrl_4;
          end
        end
        th_ctrl_3: begin
          _th_ctrl_i_0 <= _th_ctrl_i_0 + 1;
          th_ctrl <= th_ctrl_2;
        end
        th_ctrl_4: begin
          if((__saxi_outstanding_wcount == 0) && (_saxi_awready || !_saxi_awvalid)) begin
            th_ctrl <= th_ctrl_5;
          end 
        end
        th_ctrl_5: begin
          if(_saxi_awvalid && _saxi_awready) begin
            th_ctrl <= th_ctrl_6;
          end 
        end
        th_ctrl_6: begin
          if(__saxi_wready_sb_0 || !__saxi_wvalid_sb_0) begin
            th_ctrl <= th_ctrl_7;
          end 
        end
        th_ctrl_7: begin
          if(__saxi_wvalid_sb_0 && __saxi_wready_sb_0) begin
            th_ctrl <= th_ctrl_8;
          end 
        end
        th_ctrl_8: begin
          if(!__saxi_has_outstanding_write) begin
            th_ctrl <= th_ctrl_9;
          end 
        end
        th_ctrl_9: begin
          _th_ctrl_start_time_1 <= time_counter;
          th_ctrl <= th_ctrl_10;
        end
        th_ctrl_10: begin
          if((__saxi_outstanding_wcount == 0) && (_saxi_awready || !_saxi_awvalid)) begin
            th_ctrl <= th_ctrl_11;
          end 
        end
        th_ctrl_11: begin
          if(_saxi_awvalid && _saxi_awready) begin
            th_ctrl <= th_ctrl_12;
          end 
        end
        th_ctrl_12: begin
          if(__saxi_wready_sb_0 || !__saxi_wvalid_sb_0) begin
            th_ctrl <= th_ctrl_13;
          end 
        end
        th_ctrl_13: begin
          if(__saxi_wvalid_sb_0 && __saxi_wready_sb_0) begin
            th_ctrl <= th_ctrl_14;
          end 
        end
        th_ctrl_14: begin
          if(!__saxi_has_outstanding_write) begin
            th_ctrl <= th_ctrl_15;
          end 
        end
        th_ctrl_15: begin
          if(_saxi_arready || !_saxi_arvalid) begin
            th_ctrl <= th_ctrl_16;
          end 
        end
        th_ctrl_16: begin
          if(_saxi_arvalid && _saxi_arready) begin
            th_ctrl <= th_ctrl_17;
          end 
        end
        th_ctrl_17: begin
          if(__saxi_rvalid_sb_0) begin
            axim_rdata_73 <= __saxi_rdata_sb_0;
          end 
          if(__saxi_rvalid_sb_0) begin
            th_ctrl <= th_ctrl_18;
          end 
        end
        th_ctrl_18: begin
          if(axim_rdata_73 != 0) begin
            th_ctrl <= th_ctrl_15;
          end 
          if(axim_rdata_73 == 0) begin
            th_ctrl <= th_ctrl_19;
          end 
        end
        th_ctrl_19: begin
          $display("# start");
          th_ctrl <= th_ctrl_20;
        end
        th_ctrl_20: begin
          if(_saxi_arready || !_saxi_arvalid) begin
            th_ctrl <= th_ctrl_21;
          end 
        end
        th_ctrl_21: begin
          if(_saxi_arvalid && _saxi_arready) begin
            th_ctrl <= th_ctrl_22;
          end 
        end
        th_ctrl_22: begin
          if(__saxi_rvalid_sb_0) begin
            axim_rdata_74 <= __saxi_rdata_sb_0;
          end 
          if(__saxi_rvalid_sb_0) begin
            th_ctrl <= th_ctrl_23;
          end 
        end
        th_ctrl_23: begin
          if(axim_rdata_74 != 0) begin
            th_ctrl <= th_ctrl_20;
          end 
          if(axim_rdata_74 == 0) begin
            th_ctrl <= th_ctrl_24;
          end 
        end
        th_ctrl_24: begin
          _th_ctrl_end_time_2 <= time_counter;
          th_ctrl <= th_ctrl_25;
        end
        th_ctrl_25: begin
          $display("# end");
          th_ctrl <= th_ctrl_26;
        end
        th_ctrl_26: begin
          $display("# execution cycles: %d", (_th_ctrl_end_time_2 - _th_ctrl_start_time_1));
          th_ctrl <= th_ctrl_27;
        end
        th_ctrl_27: begin
          _th_ctrl_ok_3 <= 1;
          th_ctrl <= th_ctrl_28;
        end
        th_ctrl_28: begin
          _th_ctrl_bat_4 <= 0;
          th_ctrl <= th_ctrl_29;
        end
        th_ctrl_29: begin
          if(_th_ctrl_bat_4 < 1) begin
            th_ctrl <= th_ctrl_30;
          end else begin
            th_ctrl <= th_ctrl_43;
          end
        end
        th_ctrl_30: begin
          _th_ctrl_x_5 <= 0;
          th_ctrl <= th_ctrl_31;
        end
        th_ctrl_31: begin
          if(_th_ctrl_x_5 < 10) begin
            th_ctrl <= th_ctrl_32;
          end else begin
            th_ctrl <= th_ctrl_42;
          end
        end
        th_ctrl_32: begin
          if(th_ctrl == 32) begin
            rdata_75 <= { _memory_mem[0 + (_th_ctrl_bat_4 * 10 + _th_ctrl_x_5) * 16 / 8 + 1], _memory_mem[0 + (_th_ctrl_bat_4 * 10 + _th_ctrl_x_5) * 16 / 8 + 0] } >> (_th_ctrl_bat_4 * 10 + _th_ctrl_x_5) * 16 % 8;
          end 
          th_ctrl <= th_ctrl_33;
        end
        th_ctrl_33: begin
          _th_ctrl_orig_6 <= rdata_75;
          th_ctrl <= th_ctrl_34;
        end
        th_ctrl_34: begin
          if(th_ctrl == 34) begin
            rdata_76 <= { _memory_mem[8481984 + (_th_ctrl_bat_4 * 10 + _th_ctrl_x_5) * 16 / 8 + 1], _memory_mem[8481984 + (_th_ctrl_bat_4 * 10 + _th_ctrl_x_5) * 16 / 8 + 0] } >> (_th_ctrl_bat_4 * 10 + _th_ctrl_x_5) * 16 % 8;
          end 
          th_ctrl <= th_ctrl_35;
        end
        th_ctrl_35: begin
          _th_ctrl_check_7 <= rdata_76;
          th_ctrl <= th_ctrl_36;
        end
        th_ctrl_36: begin
          if(_th_ctrl_orig_6 !== _th_ctrl_check_7) begin
            th_ctrl <= th_ctrl_37;
          end else begin
            th_ctrl <= th_ctrl_40;
          end
        end
        th_ctrl_37: begin
          $display("NG ( %d %d ) orig:  %d  check:  %d", _th_ctrl_bat_4, _th_ctrl_x_5, _th_ctrl_orig_6, _th_ctrl_check_7);
          th_ctrl <= th_ctrl_38;
        end
        th_ctrl_38: begin
          _th_ctrl_ok_3 <= 0;
          th_ctrl <= th_ctrl_39;
        end
        th_ctrl_39: begin
          th_ctrl <= th_ctrl_41;
        end
        th_ctrl_40: begin
          $display("OK ( %d %d ) orig:  %d  check:  %d", _th_ctrl_bat_4, _th_ctrl_x_5, _th_ctrl_orig_6, _th_ctrl_check_7);
          th_ctrl <= th_ctrl_41;
        end
        th_ctrl_41: begin
          _th_ctrl_x_5 <= _th_ctrl_x_5 + 1;
          th_ctrl <= th_ctrl_31;
        end
        th_ctrl_42: begin
          _th_ctrl_bat_4 <= _th_ctrl_bat_4 + 1;
          th_ctrl <= th_ctrl_29;
        end
        th_ctrl_43: begin
          if(_th_ctrl_ok_3) begin
            th_ctrl <= th_ctrl_44;
          end else begin
            th_ctrl <= th_ctrl_46;
          end
        end
        th_ctrl_44: begin
          $display("# verify: PASSED");
          th_ctrl <= th_ctrl_45;
        end
        th_ctrl_45: begin
          th_ctrl <= th_ctrl_47;
        end
        th_ctrl_46: begin
          $display("# verify: FAILED");
          th_ctrl <= th_ctrl_47;
        end
        th_ctrl_47: begin
          $finish;
          th_ctrl <= th_ctrl_48;
        end
      endcase
    end
  end


endmodule



module _memory_wreq_fifo
(
  input CLK,
  input RST,
  input _memory_wreq_fifo_enq,
  input [41-1:0] _memory_wreq_fifo_wdata,
  output _memory_wreq_fifo_full,
  output _memory_wreq_fifo_almost_full,
  input _memory_wreq_fifo_deq,
  output [41-1:0] _memory_wreq_fifo_rdata,
  output _memory_wreq_fifo_empty,
  output _memory_wreq_fifo_almost_empty
);

  reg [41-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [41-1:0] rdata;
  assign _memory_wreq_fifo_full = is_full;
  assign _memory_wreq_fifo_almost_full = is_almost_full || is_full;
  assign _memory_wreq_fifo_empty = is_empty;
  assign _memory_wreq_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _memory_wreq_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_memory_wreq_fifo_enq && !is_full) begin
        mem[head] <= _memory_wreq_fifo_wdata;
        head <= head + 1;
      end 
      if(_memory_wreq_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _memory_rreq_fifo
(
  input CLK,
  input RST,
  input _memory_rreq_fifo_enq,
  input [41-1:0] _memory_rreq_fifo_wdata,
  output _memory_rreq_fifo_full,
  output _memory_rreq_fifo_almost_full,
  input _memory_rreq_fifo_deq,
  output [41-1:0] _memory_rreq_fifo_rdata,
  output _memory_rreq_fifo_empty,
  output _memory_rreq_fifo_almost_empty
);

  reg [41-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [41-1:0] rdata;
  assign _memory_rreq_fifo_full = is_full;
  assign _memory_rreq_fifo_almost_full = is_almost_full || is_full;
  assign _memory_rreq_fifo_empty = is_empty;
  assign _memory_rreq_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _memory_rreq_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_memory_rreq_fifo_enq && !is_full) begin
        mem[head] <= _memory_rreq_fifo_wdata;
        head <= head + 1;
      end 
      if(_memory_rreq_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _memory_wdata_fifo
(
  input CLK,
  input RST,
  input _memory_wdata_fifo_enq,
  input [37-1:0] _memory_wdata_fifo_wdata,
  output _memory_wdata_fifo_full,
  output _memory_wdata_fifo_almost_full,
  input _memory_wdata_fifo_deq,
  output [37-1:0] _memory_wdata_fifo_rdata,
  output _memory_wdata_fifo_empty,
  output _memory_wdata_fifo_almost_empty
);

  reg [37-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [37-1:0] rdata;
  assign _memory_wdata_fifo_full = is_full;
  assign _memory_wdata_fifo_almost_full = is_almost_full || is_full;
  assign _memory_wdata_fifo_empty = is_empty;
  assign _memory_wdata_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _memory_wdata_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_memory_wdata_fifo_enq && !is_full) begin
        mem[head] <= _memory_wdata_fifo_wdata;
        head <= head + 1;
      end 
      if(_memory_wdata_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module hello_nngen
(
  input CLK,
  input RESETN,
  output reg irq,
  output reg [32-1:0] maxi_awaddr,
  output reg [8-1:0] maxi_awlen,
  output [3-1:0] maxi_awsize,
  output [2-1:0] maxi_awburst,
  output [1-1:0] maxi_awlock,
  output [4-1:0] maxi_awcache,
  output [3-1:0] maxi_awprot,
  output [4-1:0] maxi_awqos,
  output [2-1:0] maxi_awuser,
  output reg maxi_awvalid,
  input maxi_awready,
  output [32-1:0] maxi_wdata,
  output [4-1:0] maxi_wstrb,
  output maxi_wlast,
  output maxi_wvalid,
  input maxi_wready,
  input [2-1:0] maxi_bresp,
  input maxi_bvalid,
  output maxi_bready,
  output reg [32-1:0] maxi_araddr,
  output reg [8-1:0] maxi_arlen,
  output [3-1:0] maxi_arsize,
  output [2-1:0] maxi_arburst,
  output [1-1:0] maxi_arlock,
  output [4-1:0] maxi_arcache,
  output [3-1:0] maxi_arprot,
  output [4-1:0] maxi_arqos,
  output [2-1:0] maxi_aruser,
  output reg maxi_arvalid,
  input maxi_arready,
  input [32-1:0] maxi_rdata,
  input [2-1:0] maxi_rresp,
  input maxi_rlast,
  input maxi_rvalid,
  output maxi_rready,
  input [32-1:0] saxi_awaddr,
  input [4-1:0] saxi_awcache,
  input [3-1:0] saxi_awprot,
  input saxi_awvalid,
  output saxi_awready,
  input [32-1:0] saxi_wdata,
  input [4-1:0] saxi_wstrb,
  input saxi_wvalid,
  output saxi_wready,
  output [2-1:0] saxi_bresp,
  output reg saxi_bvalid,
  input saxi_bready,
  input [32-1:0] saxi_araddr,
  input [4-1:0] saxi_arcache,
  input [3-1:0] saxi_arprot,
  input saxi_arvalid,
  output saxi_arready,
  output reg [32-1:0] saxi_rdata,
  output [2-1:0] saxi_rresp,
  output reg saxi_rvalid,
  input saxi_rready
);

  wire RESETN_inv;
  assign RESETN_inv = !RESETN;
  wire RESETN_inv_buf;
  reg _RESETN_inv_1;
  reg _RESETN_inv_2;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign maxi_awsize = 2;
  assign maxi_awburst = 1;
  assign maxi_awlock = 0;
  assign maxi_awcache = 3;
  assign maxi_awprot = 0;
  assign maxi_awqos = 0;
  assign maxi_awuser = 0;
  reg [32-1:0] _maxi_wdata_sb_0;
  reg [4-1:0] _maxi_wstrb_sb_0;
  reg _maxi_wlast_sb_0;
  reg _maxi_wvalid_sb_0;
  wire _maxi_wready_sb_0;
  wire _sb_maxi_writedata_s_value_0;
  assign _sb_maxi_writedata_s_value_0 = _maxi_wlast_sb_0;
  wire [4-1:0] _sb_maxi_writedata_s_value_1;
  assign _sb_maxi_writedata_s_value_1 = _maxi_wstrb_sb_0;
  wire [32-1:0] _sb_maxi_writedata_s_value_2;
  assign _sb_maxi_writedata_s_value_2 = _maxi_wdata_sb_0;
  wire [37-1:0] _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_s_data_3 = { _sb_maxi_writedata_s_value_0, _sb_maxi_writedata_s_value_1, _sb_maxi_writedata_s_value_2 };
  wire _sb_maxi_writedata_s_valid_4;
  assign _sb_maxi_writedata_s_valid_4 = _maxi_wvalid_sb_0;
  wire _sb_maxi_writedata_m_ready_5;
  assign _sb_maxi_writedata_m_ready_5 = maxi_wready;
  reg [37-1:0] _sb_maxi_writedata_data_6;
  reg _sb_maxi_writedata_valid_7;
  wire _sb_maxi_writedata_ready_8;
  reg [37-1:0] _sb_maxi_writedata_tmp_data_9;
  reg _sb_maxi_writedata_tmp_valid_10;
  wire [37-1:0] _sb_maxi_writedata_next_data_11;
  wire _sb_maxi_writedata_next_valid_12;
  assign _sb_maxi_writedata_ready_8 = !_sb_maxi_writedata_tmp_valid_10;
  assign _sb_maxi_writedata_next_data_11 = (_sb_maxi_writedata_tmp_valid_10)? _sb_maxi_writedata_tmp_data_9 : _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_next_valid_12 = _sb_maxi_writedata_tmp_valid_10 || _sb_maxi_writedata_s_valid_4;
  wire _sb_maxi_writedata_m_value_13;
  assign _sb_maxi_writedata_m_value_13 = _sb_maxi_writedata_data_6[36:36];
  wire [4-1:0] _sb_maxi_writedata_m_value_14;
  assign _sb_maxi_writedata_m_value_14 = _sb_maxi_writedata_data_6[35:32];
  wire [32-1:0] _sb_maxi_writedata_m_value_15;
  assign _sb_maxi_writedata_m_value_15 = _sb_maxi_writedata_data_6[31:0];
  assign _maxi_wready_sb_0 = _sb_maxi_writedata_ready_8;
  assign maxi_wdata = _sb_maxi_writedata_m_value_15;
  assign maxi_wstrb = _sb_maxi_writedata_m_value_14;
  assign maxi_wlast = _sb_maxi_writedata_m_value_13;
  assign maxi_wvalid = _sb_maxi_writedata_valid_7;
  assign maxi_bready = 1;
  assign maxi_arsize = 2;
  assign maxi_arburst = 1;
  assign maxi_arlock = 0;
  assign maxi_arcache = 3;
  assign maxi_arprot = 0;
  assign maxi_arqos = 0;
  assign maxi_aruser = 0;
  wire [32-1:0] _maxi_rdata_sb_0;
  wire _maxi_rlast_sb_0;
  wire _maxi_rvalid_sb_0;
  wire _maxi_rready_sb_0;
  wire _sb_maxi_readdata_s_value_16;
  assign _sb_maxi_readdata_s_value_16 = maxi_rlast;
  wire [32-1:0] _sb_maxi_readdata_s_value_17;
  assign _sb_maxi_readdata_s_value_17 = maxi_rdata;
  wire [33-1:0] _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_s_data_18 = { _sb_maxi_readdata_s_value_16, _sb_maxi_readdata_s_value_17 };
  wire _sb_maxi_readdata_s_valid_19;
  assign _sb_maxi_readdata_s_valid_19 = maxi_rvalid;
  wire _sb_maxi_readdata_m_ready_20;
  assign _sb_maxi_readdata_m_ready_20 = _maxi_rready_sb_0;
  reg [33-1:0] _sb_maxi_readdata_data_21;
  reg _sb_maxi_readdata_valid_22;
  wire _sb_maxi_readdata_ready_23;
  reg [33-1:0] _sb_maxi_readdata_tmp_data_24;
  reg _sb_maxi_readdata_tmp_valid_25;
  wire [33-1:0] _sb_maxi_readdata_next_data_26;
  wire _sb_maxi_readdata_next_valid_27;
  assign _sb_maxi_readdata_ready_23 = !_sb_maxi_readdata_tmp_valid_25;
  assign _sb_maxi_readdata_next_data_26 = (_sb_maxi_readdata_tmp_valid_25)? _sb_maxi_readdata_tmp_data_24 : _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_next_valid_27 = _sb_maxi_readdata_tmp_valid_25 || _sb_maxi_readdata_s_valid_19;
  wire _sb_maxi_readdata_m_value_28;
  assign _sb_maxi_readdata_m_value_28 = _sb_maxi_readdata_data_21[32:32];
  wire [32-1:0] _sb_maxi_readdata_m_value_29;
  assign _sb_maxi_readdata_m_value_29 = _sb_maxi_readdata_data_21[31:0];
  assign _maxi_rdata_sb_0 = _sb_maxi_readdata_m_value_29;
  assign _maxi_rlast_sb_0 = _sb_maxi_readdata_m_value_28;
  assign _maxi_rvalid_sb_0 = _sb_maxi_readdata_valid_22;
  assign maxi_rready = _sb_maxi_readdata_ready_23;
  reg [3-1:0] _maxi_outstanding_wcount;
  wire _maxi_has_outstanding_write;
  assign _maxi_has_outstanding_write = (_maxi_outstanding_wcount > 0) || maxi_awvalid;
  reg _maxi_read_start;
  reg [8-1:0] _maxi_read_op_sel;
  reg [32-1:0] _maxi_read_global_addr;
  reg [33-1:0] _maxi_read_global_size;
  reg [32-1:0] _maxi_read_local_addr;
  reg [32-1:0] _maxi_read_local_stride;
  reg [33-1:0] _maxi_read_local_size;
  reg [32-1:0] _maxi_read_local_blocksize;
  wire _maxi_read_req_fifo_enq;
  wire [137-1:0] _maxi_read_req_fifo_wdata;
  wire _maxi_read_req_fifo_full;
  wire _maxi_read_req_fifo_almost_full;
  wire _maxi_read_req_fifo_deq;
  wire [137-1:0] _maxi_read_req_fifo_rdata;
  wire _maxi_read_req_fifo_empty;
  wire _maxi_read_req_fifo_almost_empty;

  _maxi_read_req_fifo
  inst__maxi_read_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_read_req_fifo_enq(_maxi_read_req_fifo_enq),
    ._maxi_read_req_fifo_wdata(_maxi_read_req_fifo_wdata),
    ._maxi_read_req_fifo_full(_maxi_read_req_fifo_full),
    ._maxi_read_req_fifo_almost_full(_maxi_read_req_fifo_almost_full),
    ._maxi_read_req_fifo_deq(_maxi_read_req_fifo_deq),
    ._maxi_read_req_fifo_rdata(_maxi_read_req_fifo_rdata),
    ._maxi_read_req_fifo_empty(_maxi_read_req_fifo_empty),
    ._maxi_read_req_fifo_almost_empty(_maxi_read_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_read_req_fifo;
  wire [8-1:0] _maxi_read_op_sel_fifo;
  wire [32-1:0] _maxi_read_local_addr_fifo;
  wire [32-1:0] _maxi_read_local_stride_fifo;
  wire [33-1:0] _maxi_read_local_size_fifo;
  wire [32-1:0] _maxi_read_local_blocksize_fifo;
  wire [8-1:0] unpack_read_req_op_sel_30;
  wire [32-1:0] unpack_read_req_local_addr_31;
  wire [32-1:0] unpack_read_req_local_stride_32;
  wire [33-1:0] unpack_read_req_local_size_33;
  wire [32-1:0] unpack_read_req_local_blocksize_34;
  assign unpack_read_req_op_sel_30 = _maxi_read_req_fifo_rdata[136:129];
  assign unpack_read_req_local_addr_31 = _maxi_read_req_fifo_rdata[128:97];
  assign unpack_read_req_local_stride_32 = _maxi_read_req_fifo_rdata[96:65];
  assign unpack_read_req_local_size_33 = _maxi_read_req_fifo_rdata[64:32];
  assign unpack_read_req_local_blocksize_34 = _maxi_read_req_fifo_rdata[31:0];
  assign _maxi_read_op_sel_fifo = unpack_read_req_op_sel_30;
  assign _maxi_read_local_addr_fifo = unpack_read_req_local_addr_31;
  assign _maxi_read_local_stride_fifo = unpack_read_req_local_stride_32;
  assign _maxi_read_local_size_fifo = unpack_read_req_local_size_33;
  assign _maxi_read_local_blocksize_fifo = unpack_read_req_local_blocksize_34;
  reg [8-1:0] _maxi_read_op_sel_buf;
  reg [32-1:0] _maxi_read_local_addr_buf;
  reg [32-1:0] _maxi_read_local_stride_buf;
  reg [33-1:0] _maxi_read_local_size_buf;
  reg [32-1:0] _maxi_read_local_blocksize_buf;
  reg _maxi_read_req_busy;
  reg _maxi_read_data_busy;
  wire _maxi_read_req_idle;
  wire _maxi_read_data_idle;
  wire _maxi_read_idle;
  assign _maxi_read_req_idle = !_maxi_read_start && !_maxi_read_req_busy;
  assign _maxi_read_data_idle = _maxi_read_req_fifo_empty && !_maxi_read_data_busy;
  assign _maxi_read_idle = _maxi_read_req_idle && _maxi_read_data_idle;
  reg _maxi_write_start;
  reg [8-1:0] _maxi_write_op_sel;
  reg [32-1:0] _maxi_write_global_addr;
  reg [33-1:0] _maxi_write_global_size;
  reg [32-1:0] _maxi_write_local_addr;
  reg [32-1:0] _maxi_write_local_stride;
  reg [33-1:0] _maxi_write_local_size;
  reg [32-1:0] _maxi_write_local_blocksize;
  wire _maxi_write_req_fifo_enq;
  wire [137-1:0] _maxi_write_req_fifo_wdata;
  wire _maxi_write_req_fifo_full;
  wire _maxi_write_req_fifo_almost_full;
  wire _maxi_write_req_fifo_deq;
  wire [137-1:0] _maxi_write_req_fifo_rdata;
  wire _maxi_write_req_fifo_empty;
  wire _maxi_write_req_fifo_almost_empty;

  _maxi_write_req_fifo
  inst__maxi_write_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_write_req_fifo_enq(_maxi_write_req_fifo_enq),
    ._maxi_write_req_fifo_wdata(_maxi_write_req_fifo_wdata),
    ._maxi_write_req_fifo_full(_maxi_write_req_fifo_full),
    ._maxi_write_req_fifo_almost_full(_maxi_write_req_fifo_almost_full),
    ._maxi_write_req_fifo_deq(_maxi_write_req_fifo_deq),
    ._maxi_write_req_fifo_rdata(_maxi_write_req_fifo_rdata),
    ._maxi_write_req_fifo_empty(_maxi_write_req_fifo_empty),
    ._maxi_write_req_fifo_almost_empty(_maxi_write_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_write_req_fifo;
  wire [8-1:0] _maxi_write_op_sel_fifo;
  wire [32-1:0] _maxi_write_local_addr_fifo;
  wire [32-1:0] _maxi_write_local_stride_fifo;
  wire [33-1:0] _maxi_write_size_fifo;
  wire [32-1:0] _maxi_write_local_blocksize_fifo;
  wire [8-1:0] unpack_write_req_op_sel_35;
  wire [32-1:0] unpack_write_req_local_addr_36;
  wire [32-1:0] unpack_write_req_local_stride_37;
  wire [33-1:0] unpack_write_req_size_38;
  wire [32-1:0] unpack_write_req_local_blocksize_39;
  assign unpack_write_req_op_sel_35 = _maxi_write_req_fifo_rdata[136:129];
  assign unpack_write_req_local_addr_36 = _maxi_write_req_fifo_rdata[128:97];
  assign unpack_write_req_local_stride_37 = _maxi_write_req_fifo_rdata[96:65];
  assign unpack_write_req_size_38 = _maxi_write_req_fifo_rdata[64:32];
  assign unpack_write_req_local_blocksize_39 = _maxi_write_req_fifo_rdata[31:0];
  assign _maxi_write_op_sel_fifo = unpack_write_req_op_sel_35;
  assign _maxi_write_local_addr_fifo = unpack_write_req_local_addr_36;
  assign _maxi_write_local_stride_fifo = unpack_write_req_local_stride_37;
  assign _maxi_write_size_fifo = unpack_write_req_size_38;
  assign _maxi_write_local_blocksize_fifo = unpack_write_req_local_blocksize_39;
  reg [8-1:0] _maxi_write_op_sel_buf;
  reg [32-1:0] _maxi_write_local_addr_buf;
  reg [32-1:0] _maxi_write_local_stride_buf;
  reg [33-1:0] _maxi_write_size_buf;
  reg [32-1:0] _maxi_write_local_blocksize_buf;
  reg _maxi_write_req_busy;
  reg _maxi_write_data_busy;
  wire _maxi_write_req_idle;
  wire _maxi_write_data_idle;
  wire _maxi_write_idle;
  assign _maxi_write_req_idle = !_maxi_write_start && !_maxi_write_req_busy;
  assign _maxi_write_data_idle = _maxi_write_req_fifo_empty && !_maxi_write_data_busy;
  assign _maxi_write_idle = _maxi_write_req_idle && _maxi_write_data_idle;
  reg [32-1:0] _maxi_global_base_addr;
  assign saxi_bresp = 0;
  assign saxi_rresp = 0;
  reg signed [32-1:0] _saxi_register_0;
  reg signed [32-1:0] _saxi_register_1;
  reg signed [32-1:0] _saxi_register_2;
  reg signed [32-1:0] _saxi_register_3;
  reg signed [32-1:0] _saxi_register_4;
  reg signed [32-1:0] _saxi_register_5;
  reg signed [32-1:0] _saxi_register_6;
  reg signed [32-1:0] _saxi_register_7;
  reg signed [32-1:0] _saxi_register_8;
  reg signed [32-1:0] _saxi_register_9;
  reg signed [32-1:0] _saxi_register_10;
  reg signed [32-1:0] _saxi_register_11;
  reg signed [32-1:0] _saxi_register_12;
  reg signed [32-1:0] _saxi_register_13;
  reg signed [32-1:0] _saxi_register_14;
  reg signed [32-1:0] _saxi_register_15;
  reg signed [32-1:0] _saxi_register_16;
  reg signed [32-1:0] _saxi_register_17;
  reg signed [32-1:0] _saxi_register_18;
  reg signed [32-1:0] _saxi_register_19;
  reg signed [32-1:0] _saxi_register_20;
  reg signed [32-1:0] _saxi_register_21;
  reg signed [32-1:0] _saxi_register_22;
  reg signed [32-1:0] _saxi_register_23;
  reg signed [32-1:0] _saxi_register_24;
  reg signed [32-1:0] _saxi_register_25;
  reg signed [32-1:0] _saxi_register_26;
  reg signed [32-1:0] _saxi_register_27;
  reg signed [32-1:0] _saxi_register_28;
  reg signed [32-1:0] _saxi_register_29;
  reg signed [32-1:0] _saxi_register_30;
  reg signed [32-1:0] _saxi_register_31;
  reg signed [32-1:0] _saxi_register_32;
  reg signed [32-1:0] _saxi_register_33;
  reg signed [32-1:0] _saxi_register_34;
  reg signed [32-1:0] _saxi_register_35;
  reg signed [32-1:0] _saxi_register_36;
  reg _saxi_flag_0;
  reg _saxi_flag_1;
  reg _saxi_flag_2;
  reg _saxi_flag_3;
  reg _saxi_flag_4;
  reg _saxi_flag_5;
  reg _saxi_flag_6;
  reg _saxi_flag_7;
  reg _saxi_flag_8;
  reg _saxi_flag_9;
  reg _saxi_flag_10;
  reg _saxi_flag_11;
  reg _saxi_flag_12;
  reg _saxi_flag_13;
  reg _saxi_flag_14;
  reg _saxi_flag_15;
  reg _saxi_flag_16;
  reg _saxi_flag_17;
  reg _saxi_flag_18;
  reg _saxi_flag_19;
  reg _saxi_flag_20;
  reg _saxi_flag_21;
  reg _saxi_flag_22;
  reg _saxi_flag_23;
  reg _saxi_flag_24;
  reg _saxi_flag_25;
  reg _saxi_flag_26;
  reg _saxi_flag_27;
  reg _saxi_flag_28;
  reg _saxi_flag_29;
  reg _saxi_flag_30;
  reg _saxi_flag_31;
  reg _saxi_flag_32;
  reg _saxi_flag_33;
  reg _saxi_flag_34;
  reg _saxi_flag_35;
  reg _saxi_flag_36;
  reg signed [32-1:0] _saxi_resetval_0;
  reg signed [32-1:0] _saxi_resetval_1;
  reg signed [32-1:0] _saxi_resetval_2;
  reg signed [32-1:0] _saxi_resetval_3;
  reg signed [32-1:0] _saxi_resetval_4;
  reg signed [32-1:0] _saxi_resetval_5;
  reg signed [32-1:0] _saxi_resetval_6;
  reg signed [32-1:0] _saxi_resetval_7;
  reg signed [32-1:0] _saxi_resetval_8;
  reg signed [32-1:0] _saxi_resetval_9;
  reg signed [32-1:0] _saxi_resetval_10;
  reg signed [32-1:0] _saxi_resetval_11;
  reg signed [32-1:0] _saxi_resetval_12;
  reg signed [32-1:0] _saxi_resetval_13;
  reg signed [32-1:0] _saxi_resetval_14;
  reg signed [32-1:0] _saxi_resetval_15;
  reg signed [32-1:0] _saxi_resetval_16;
  reg signed [32-1:0] _saxi_resetval_17;
  reg signed [32-1:0] _saxi_resetval_18;
  reg signed [32-1:0] _saxi_resetval_19;
  reg signed [32-1:0] _saxi_resetval_20;
  reg signed [32-1:0] _saxi_resetval_21;
  reg signed [32-1:0] _saxi_resetval_22;
  reg signed [32-1:0] _saxi_resetval_23;
  reg signed [32-1:0] _saxi_resetval_24;
  reg signed [32-1:0] _saxi_resetval_25;
  reg signed [32-1:0] _saxi_resetval_26;
  reg signed [32-1:0] _saxi_resetval_27;
  reg signed [32-1:0] _saxi_resetval_28;
  reg signed [32-1:0] _saxi_resetval_29;
  reg signed [32-1:0] _saxi_resetval_30;
  reg signed [32-1:0] _saxi_resetval_31;
  reg signed [32-1:0] _saxi_resetval_32;
  reg signed [32-1:0] _saxi_resetval_33;
  reg signed [32-1:0] _saxi_resetval_34;
  reg signed [32-1:0] _saxi_resetval_35;
  reg signed [32-1:0] _saxi_resetval_36;
  localparam _saxi_maskwidth = 6;
  localparam _saxi_mask = { _saxi_maskwidth{ 1'd1 } };
  localparam _saxi_shift = 2;
  reg [32-1:0] _saxi_register_fsm;
  localparam _saxi_register_fsm_init = 0;
  reg [32-1:0] addr_40;
  reg writevalid_41;
  reg readvalid_42;
  reg prev_awvalid_43;
  reg prev_arvalid_44;
  assign saxi_awready = (_saxi_register_fsm == 0) && (!writevalid_41 && !readvalid_42 && !saxi_bvalid && prev_awvalid_43);
  assign saxi_arready = (_saxi_register_fsm == 0) && (!readvalid_42 && !writevalid_41 && prev_arvalid_44 && !prev_awvalid_43);
  reg [_saxi_maskwidth-1:0] axis_maskaddr_45;
  wire signed [32-1:0] axislite_rdata_46;
  assign axislite_rdata_46 = (axis_maskaddr_45 == 0)? _saxi_register_0 : 
                             (axis_maskaddr_45 == 1)? _saxi_register_1 : 
                             (axis_maskaddr_45 == 2)? _saxi_register_2 : 
                             (axis_maskaddr_45 == 3)? _saxi_register_3 : 
                             (axis_maskaddr_45 == 4)? _saxi_register_4 : 
                             (axis_maskaddr_45 == 5)? _saxi_register_5 : 
                             (axis_maskaddr_45 == 6)? _saxi_register_6 : 
                             (axis_maskaddr_45 == 7)? _saxi_register_7 : 
                             (axis_maskaddr_45 == 8)? _saxi_register_8 : 
                             (axis_maskaddr_45 == 9)? _saxi_register_9 : 
                             (axis_maskaddr_45 == 10)? _saxi_register_10 : 
                             (axis_maskaddr_45 == 11)? _saxi_register_11 : 
                             (axis_maskaddr_45 == 12)? _saxi_register_12 : 
                             (axis_maskaddr_45 == 13)? _saxi_register_13 : 
                             (axis_maskaddr_45 == 14)? _saxi_register_14 : 
                             (axis_maskaddr_45 == 15)? _saxi_register_15 : 
                             (axis_maskaddr_45 == 16)? _saxi_register_16 : 
                             (axis_maskaddr_45 == 17)? _saxi_register_17 : 
                             (axis_maskaddr_45 == 18)? _saxi_register_18 : 
                             (axis_maskaddr_45 == 19)? _saxi_register_19 : 
                             (axis_maskaddr_45 == 20)? _saxi_register_20 : 
                             (axis_maskaddr_45 == 21)? _saxi_register_21 : 
                             (axis_maskaddr_45 == 22)? _saxi_register_22 : 
                             (axis_maskaddr_45 == 23)? _saxi_register_23 : 
                             (axis_maskaddr_45 == 24)? _saxi_register_24 : 
                             (axis_maskaddr_45 == 25)? _saxi_register_25 : 
                             (axis_maskaddr_45 == 26)? _saxi_register_26 : 
                             (axis_maskaddr_45 == 27)? _saxi_register_27 : 
                             (axis_maskaddr_45 == 28)? _saxi_register_28 : 
                             (axis_maskaddr_45 == 29)? _saxi_register_29 : 
                             (axis_maskaddr_45 == 30)? _saxi_register_30 : 
                             (axis_maskaddr_45 == 31)? _saxi_register_31 : 
                             (axis_maskaddr_45 == 32)? _saxi_register_32 : 
                             (axis_maskaddr_45 == 33)? _saxi_register_33 : 
                             (axis_maskaddr_45 == 34)? _saxi_register_34 : 
                             (axis_maskaddr_45 == 35)? _saxi_register_35 : 
                             (axis_maskaddr_45 == 36)? _saxi_register_36 : 'hx;
  wire axislite_flag_47;
  assign axislite_flag_47 = (axis_maskaddr_45 == 0)? _saxi_flag_0 : 
                            (axis_maskaddr_45 == 1)? _saxi_flag_1 : 
                            (axis_maskaddr_45 == 2)? _saxi_flag_2 : 
                            (axis_maskaddr_45 == 3)? _saxi_flag_3 : 
                            (axis_maskaddr_45 == 4)? _saxi_flag_4 : 
                            (axis_maskaddr_45 == 5)? _saxi_flag_5 : 
                            (axis_maskaddr_45 == 6)? _saxi_flag_6 : 
                            (axis_maskaddr_45 == 7)? _saxi_flag_7 : 
                            (axis_maskaddr_45 == 8)? _saxi_flag_8 : 
                            (axis_maskaddr_45 == 9)? _saxi_flag_9 : 
                            (axis_maskaddr_45 == 10)? _saxi_flag_10 : 
                            (axis_maskaddr_45 == 11)? _saxi_flag_11 : 
                            (axis_maskaddr_45 == 12)? _saxi_flag_12 : 
                            (axis_maskaddr_45 == 13)? _saxi_flag_13 : 
                            (axis_maskaddr_45 == 14)? _saxi_flag_14 : 
                            (axis_maskaddr_45 == 15)? _saxi_flag_15 : 
                            (axis_maskaddr_45 == 16)? _saxi_flag_16 : 
                            (axis_maskaddr_45 == 17)? _saxi_flag_17 : 
                            (axis_maskaddr_45 == 18)? _saxi_flag_18 : 
                            (axis_maskaddr_45 == 19)? _saxi_flag_19 : 
                            (axis_maskaddr_45 == 20)? _saxi_flag_20 : 
                            (axis_maskaddr_45 == 21)? _saxi_flag_21 : 
                            (axis_maskaddr_45 == 22)? _saxi_flag_22 : 
                            (axis_maskaddr_45 == 23)? _saxi_flag_23 : 
                            (axis_maskaddr_45 == 24)? _saxi_flag_24 : 
                            (axis_maskaddr_45 == 25)? _saxi_flag_25 : 
                            (axis_maskaddr_45 == 26)? _saxi_flag_26 : 
                            (axis_maskaddr_45 == 27)? _saxi_flag_27 : 
                            (axis_maskaddr_45 == 28)? _saxi_flag_28 : 
                            (axis_maskaddr_45 == 29)? _saxi_flag_29 : 
                            (axis_maskaddr_45 == 30)? _saxi_flag_30 : 
                            (axis_maskaddr_45 == 31)? _saxi_flag_31 : 
                            (axis_maskaddr_45 == 32)? _saxi_flag_32 : 
                            (axis_maskaddr_45 == 33)? _saxi_flag_33 : 
                            (axis_maskaddr_45 == 34)? _saxi_flag_34 : 
                            (axis_maskaddr_45 == 35)? _saxi_flag_35 : 
                            (axis_maskaddr_45 == 36)? _saxi_flag_36 : 'hx;
  wire signed [32-1:0] axislite_resetval_48;
  assign axislite_resetval_48 = (axis_maskaddr_45 == 0)? _saxi_resetval_0 : 
                                (axis_maskaddr_45 == 1)? _saxi_resetval_1 : 
                                (axis_maskaddr_45 == 2)? _saxi_resetval_2 : 
                                (axis_maskaddr_45 == 3)? _saxi_resetval_3 : 
                                (axis_maskaddr_45 == 4)? _saxi_resetval_4 : 
                                (axis_maskaddr_45 == 5)? _saxi_resetval_5 : 
                                (axis_maskaddr_45 == 6)? _saxi_resetval_6 : 
                                (axis_maskaddr_45 == 7)? _saxi_resetval_7 : 
                                (axis_maskaddr_45 == 8)? _saxi_resetval_8 : 
                                (axis_maskaddr_45 == 9)? _saxi_resetval_9 : 
                                (axis_maskaddr_45 == 10)? _saxi_resetval_10 : 
                                (axis_maskaddr_45 == 11)? _saxi_resetval_11 : 
                                (axis_maskaddr_45 == 12)? _saxi_resetval_12 : 
                                (axis_maskaddr_45 == 13)? _saxi_resetval_13 : 
                                (axis_maskaddr_45 == 14)? _saxi_resetval_14 : 
                                (axis_maskaddr_45 == 15)? _saxi_resetval_15 : 
                                (axis_maskaddr_45 == 16)? _saxi_resetval_16 : 
                                (axis_maskaddr_45 == 17)? _saxi_resetval_17 : 
                                (axis_maskaddr_45 == 18)? _saxi_resetval_18 : 
                                (axis_maskaddr_45 == 19)? _saxi_resetval_19 : 
                                (axis_maskaddr_45 == 20)? _saxi_resetval_20 : 
                                (axis_maskaddr_45 == 21)? _saxi_resetval_21 : 
                                (axis_maskaddr_45 == 22)? _saxi_resetval_22 : 
                                (axis_maskaddr_45 == 23)? _saxi_resetval_23 : 
                                (axis_maskaddr_45 == 24)? _saxi_resetval_24 : 
                                (axis_maskaddr_45 == 25)? _saxi_resetval_25 : 
                                (axis_maskaddr_45 == 26)? _saxi_resetval_26 : 
                                (axis_maskaddr_45 == 27)? _saxi_resetval_27 : 
                                (axis_maskaddr_45 == 28)? _saxi_resetval_28 : 
                                (axis_maskaddr_45 == 29)? _saxi_resetval_29 : 
                                (axis_maskaddr_45 == 30)? _saxi_resetval_30 : 
                                (axis_maskaddr_45 == 31)? _saxi_resetval_31 : 
                                (axis_maskaddr_45 == 32)? _saxi_resetval_32 : 
                                (axis_maskaddr_45 == 33)? _saxi_resetval_33 : 
                                (axis_maskaddr_45 == 34)? _saxi_resetval_34 : 
                                (axis_maskaddr_45 == 35)? _saxi_resetval_35 : 
                                (axis_maskaddr_45 == 36)? _saxi_resetval_36 : 'hx;
  reg _saxi_rdata_cond_0_1;
  assign saxi_wready = _saxi_register_fsm == 3;
  wire maxi_idle;
  assign maxi_idle = _maxi_write_idle & _maxi_read_idle;
  wire sw_rst_logic;
  assign sw_rst_logic = maxi_idle & _saxi_register_6;
  wire rst_logic;
  assign rst_logic = RESETN_inv_buf | sw_rst_logic;
  reg RST;
  reg _rst_logic_1;
  reg _rst_logic_2;
  wire signed [32-1:0] irq_49;
  assign irq_49 = _saxi_register_9 & _saxi_register_10;
  wire irq_busy;
  assign irq_busy = _saxi_register_5[0];
  reg irq_busy_edge_50;
  wire irq_busy_edge_51;
  assign irq_busy_edge_51 = irq_busy_edge_50 & !irq_busy;
  wire irq_extern;
  assign irq_extern = |_saxi_register_7;
  reg irq_extern_edge_52;
  wire irq_extern_edge_53;
  assign irq_extern_edge_53 = !irq_extern_edge_52 & irq_extern;
  wire [14-1:0] ram_w32_l16384_id0_0_addr;
  wire [32-1:0] ram_w32_l16384_id0_0_rdata;
  wire [32-1:0] ram_w32_l16384_id0_0_wdata;
  wire ram_w32_l16384_id0_0_wenable;
  wire ram_w32_l16384_id0_0_enable;
  wire [14-1:0] ram_w32_l16384_id0_1_addr;
  wire [32-1:0] ram_w32_l16384_id0_1_rdata;
  wire [32-1:0] ram_w32_l16384_id0_1_wdata;
  wire ram_w32_l16384_id0_1_wenable;
  wire ram_w32_l16384_id0_1_enable;
  assign ram_w32_l16384_id0_0_wdata = 'hx;
  assign ram_w32_l16384_id0_0_wenable = 0;

  ram_w32_l16384_id0
  inst_ram_w32_l16384_id0
  (
    .CLK(CLK),
    .ram_w32_l16384_id0_0_addr(ram_w32_l16384_id0_0_addr),
    .ram_w32_l16384_id0_0_rdata(ram_w32_l16384_id0_0_rdata),
    .ram_w32_l16384_id0_0_wdata(ram_w32_l16384_id0_0_wdata),
    .ram_w32_l16384_id0_0_wenable(ram_w32_l16384_id0_0_wenable),
    .ram_w32_l16384_id0_0_enable(ram_w32_l16384_id0_0_enable),
    .ram_w32_l16384_id0_1_addr(ram_w32_l16384_id0_1_addr),
    .ram_w32_l16384_id0_1_rdata(ram_w32_l16384_id0_1_rdata),
    .ram_w32_l16384_id0_1_wdata(ram_w32_l16384_id0_1_wdata),
    .ram_w32_l16384_id0_1_wenable(ram_w32_l16384_id0_1_wenable),
    .ram_w32_l16384_id0_1_enable(ram_w32_l16384_id0_1_enable)
  );

  wire [14-1:0] ram_w32_l16384_id1_0_addr;
  wire [32-1:0] ram_w32_l16384_id1_0_rdata;
  wire [32-1:0] ram_w32_l16384_id1_0_wdata;
  wire ram_w32_l16384_id1_0_wenable;
  wire ram_w32_l16384_id1_0_enable;
  wire [14-1:0] ram_w32_l16384_id1_1_addr;
  wire [32-1:0] ram_w32_l16384_id1_1_rdata;
  wire [32-1:0] ram_w32_l16384_id1_1_wdata;
  wire ram_w32_l16384_id1_1_wenable;
  wire ram_w32_l16384_id1_1_enable;
  assign ram_w32_l16384_id1_0_wdata = 'hx;
  assign ram_w32_l16384_id1_0_wenable = 0;

  ram_w32_l16384_id1
  inst_ram_w32_l16384_id1
  (
    .CLK(CLK),
    .ram_w32_l16384_id1_0_addr(ram_w32_l16384_id1_0_addr),
    .ram_w32_l16384_id1_0_rdata(ram_w32_l16384_id1_0_rdata),
    .ram_w32_l16384_id1_0_wdata(ram_w32_l16384_id1_0_wdata),
    .ram_w32_l16384_id1_0_wenable(ram_w32_l16384_id1_0_wenable),
    .ram_w32_l16384_id1_0_enable(ram_w32_l16384_id1_0_enable),
    .ram_w32_l16384_id1_1_addr(ram_w32_l16384_id1_1_addr),
    .ram_w32_l16384_id1_1_rdata(ram_w32_l16384_id1_1_rdata),
    .ram_w32_l16384_id1_1_wdata(ram_w32_l16384_id1_1_wdata),
    .ram_w32_l16384_id1_1_wenable(ram_w32_l16384_id1_1_wenable),
    .ram_w32_l16384_id1_1_enable(ram_w32_l16384_id1_1_enable)
  );

  wire [13-1:0] ram_w32_l8192_id0_0_addr;
  wire [32-1:0] ram_w32_l8192_id0_0_rdata;
  wire [32-1:0] ram_w32_l8192_id0_0_wdata;
  wire ram_w32_l8192_id0_0_wenable;
  wire ram_w32_l8192_id0_0_enable;
  wire [13-1:0] ram_w32_l8192_id0_1_addr;
  wire [32-1:0] ram_w32_l8192_id0_1_rdata;
  wire [32-1:0] ram_w32_l8192_id0_1_wdata;
  wire ram_w32_l8192_id0_1_wenable;
  wire ram_w32_l8192_id0_1_enable;

  ram_w32_l8192_id0
  inst_ram_w32_l8192_id0
  (
    .CLK(CLK),
    .ram_w32_l8192_id0_0_addr(ram_w32_l8192_id0_0_addr),
    .ram_w32_l8192_id0_0_rdata(ram_w32_l8192_id0_0_rdata),
    .ram_w32_l8192_id0_0_wdata(ram_w32_l8192_id0_0_wdata),
    .ram_w32_l8192_id0_0_wenable(ram_w32_l8192_id0_0_wenable),
    .ram_w32_l8192_id0_0_enable(ram_w32_l8192_id0_0_enable),
    .ram_w32_l8192_id0_1_addr(ram_w32_l8192_id0_1_addr),
    .ram_w32_l8192_id0_1_rdata(ram_w32_l8192_id0_1_rdata),
    .ram_w32_l8192_id0_1_wdata(ram_w32_l8192_id0_1_wdata),
    .ram_w32_l8192_id0_1_wenable(ram_w32_l8192_id0_1_wenable),
    .ram_w32_l8192_id0_1_enable(ram_w32_l8192_id0_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id0_0_addr;
  wire [32-1:0] ram_w32_l512_id0_0_rdata;
  wire [32-1:0] ram_w32_l512_id0_0_wdata;
  wire ram_w32_l512_id0_0_wenable;
  wire ram_w32_l512_id0_0_enable;
  wire [9-1:0] ram_w32_l512_id0_1_addr;
  wire [32-1:0] ram_w32_l512_id0_1_rdata;
  wire [32-1:0] ram_w32_l512_id0_1_wdata;
  wire ram_w32_l512_id0_1_wenable;
  wire ram_w32_l512_id0_1_enable;
  assign ram_w32_l512_id0_0_wdata = 'hx;
  assign ram_w32_l512_id0_0_wenable = 0;

  ram_w32_l512_id0
  inst_ram_w32_l512_id0
  (
    .CLK(CLK),
    .ram_w32_l512_id0_0_addr(ram_w32_l512_id0_0_addr),
    .ram_w32_l512_id0_0_rdata(ram_w32_l512_id0_0_rdata),
    .ram_w32_l512_id0_0_wdata(ram_w32_l512_id0_0_wdata),
    .ram_w32_l512_id0_0_wenable(ram_w32_l512_id0_0_wenable),
    .ram_w32_l512_id0_0_enable(ram_w32_l512_id0_0_enable),
    .ram_w32_l512_id0_1_addr(ram_w32_l512_id0_1_addr),
    .ram_w32_l512_id0_1_rdata(ram_w32_l512_id0_1_rdata),
    .ram_w32_l512_id0_1_wdata(ram_w32_l512_id0_1_wdata),
    .ram_w32_l512_id0_1_wenable(ram_w32_l512_id0_1_wenable),
    .ram_w32_l512_id0_1_enable(ram_w32_l512_id0_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id1_0_addr;
  wire [32-1:0] ram_w32_l512_id1_0_rdata;
  wire [32-1:0] ram_w32_l512_id1_0_wdata;
  wire ram_w32_l512_id1_0_wenable;
  wire ram_w32_l512_id1_0_enable;
  wire [9-1:0] ram_w32_l512_id1_1_addr;
  wire [32-1:0] ram_w32_l512_id1_1_rdata;
  wire [32-1:0] ram_w32_l512_id1_1_wdata;
  wire ram_w32_l512_id1_1_wenable;
  wire ram_w32_l512_id1_1_enable;
  assign ram_w32_l512_id1_0_wdata = 'hx;
  assign ram_w32_l512_id1_0_wenable = 0;

  ram_w32_l512_id1
  inst_ram_w32_l512_id1
  (
    .CLK(CLK),
    .ram_w32_l512_id1_0_addr(ram_w32_l512_id1_0_addr),
    .ram_w32_l512_id1_0_rdata(ram_w32_l512_id1_0_rdata),
    .ram_w32_l512_id1_0_wdata(ram_w32_l512_id1_0_wdata),
    .ram_w32_l512_id1_0_wenable(ram_w32_l512_id1_0_wenable),
    .ram_w32_l512_id1_0_enable(ram_w32_l512_id1_0_enable),
    .ram_w32_l512_id1_1_addr(ram_w32_l512_id1_1_addr),
    .ram_w32_l512_id1_1_rdata(ram_w32_l512_id1_1_rdata),
    .ram_w32_l512_id1_1_wdata(ram_w32_l512_id1_1_wdata),
    .ram_w32_l512_id1_1_wenable(ram_w32_l512_id1_1_wenable),
    .ram_w32_l512_id1_1_enable(ram_w32_l512_id1_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id2_0_addr;
  wire [32-1:0] ram_w32_l512_id2_0_rdata;
  wire [32-1:0] ram_w32_l512_id2_0_wdata;
  wire ram_w32_l512_id2_0_wenable;
  wire ram_w32_l512_id2_0_enable;
  wire [9-1:0] ram_w32_l512_id2_1_addr;
  wire [32-1:0] ram_w32_l512_id2_1_rdata;
  wire [32-1:0] ram_w32_l512_id2_1_wdata;
  wire ram_w32_l512_id2_1_wenable;
  wire ram_w32_l512_id2_1_enable;
  assign ram_w32_l512_id2_0_wdata = 'hx;
  assign ram_w32_l512_id2_0_wenable = 0;

  ram_w32_l512_id2
  inst_ram_w32_l512_id2
  (
    .CLK(CLK),
    .ram_w32_l512_id2_0_addr(ram_w32_l512_id2_0_addr),
    .ram_w32_l512_id2_0_rdata(ram_w32_l512_id2_0_rdata),
    .ram_w32_l512_id2_0_wdata(ram_w32_l512_id2_0_wdata),
    .ram_w32_l512_id2_0_wenable(ram_w32_l512_id2_0_wenable),
    .ram_w32_l512_id2_0_enable(ram_w32_l512_id2_0_enable),
    .ram_w32_l512_id2_1_addr(ram_w32_l512_id2_1_addr),
    .ram_w32_l512_id2_1_rdata(ram_w32_l512_id2_1_rdata),
    .ram_w32_l512_id2_1_wdata(ram_w32_l512_id2_1_wdata),
    .ram_w32_l512_id2_1_wenable(ram_w32_l512_id2_1_wenable),
    .ram_w32_l512_id2_1_enable(ram_w32_l512_id2_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id3_0_addr;
  wire [32-1:0] ram_w32_l512_id3_0_rdata;
  wire [32-1:0] ram_w32_l512_id3_0_wdata;
  wire ram_w32_l512_id3_0_wenable;
  wire ram_w32_l512_id3_0_enable;
  wire [9-1:0] ram_w32_l512_id3_1_addr;
  wire [32-1:0] ram_w32_l512_id3_1_rdata;
  wire [32-1:0] ram_w32_l512_id3_1_wdata;
  wire ram_w32_l512_id3_1_wenable;
  wire ram_w32_l512_id3_1_enable;
  assign ram_w32_l512_id3_0_wdata = 'hx;
  assign ram_w32_l512_id3_0_wenable = 0;

  ram_w32_l512_id3
  inst_ram_w32_l512_id3
  (
    .CLK(CLK),
    .ram_w32_l512_id3_0_addr(ram_w32_l512_id3_0_addr),
    .ram_w32_l512_id3_0_rdata(ram_w32_l512_id3_0_rdata),
    .ram_w32_l512_id3_0_wdata(ram_w32_l512_id3_0_wdata),
    .ram_w32_l512_id3_0_wenable(ram_w32_l512_id3_0_wenable),
    .ram_w32_l512_id3_0_enable(ram_w32_l512_id3_0_enable),
    .ram_w32_l512_id3_1_addr(ram_w32_l512_id3_1_addr),
    .ram_w32_l512_id3_1_rdata(ram_w32_l512_id3_1_rdata),
    .ram_w32_l512_id3_1_wdata(ram_w32_l512_id3_1_wdata),
    .ram_w32_l512_id3_1_wenable(ram_w32_l512_id3_1_wenable),
    .ram_w32_l512_id3_1_enable(ram_w32_l512_id3_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id4_0_addr;
  wire [32-1:0] ram_w32_l512_id4_0_rdata;
  wire [32-1:0] ram_w32_l512_id4_0_wdata;
  wire ram_w32_l512_id4_0_wenable;
  wire ram_w32_l512_id4_0_enable;
  wire [9-1:0] ram_w32_l512_id4_1_addr;
  wire [32-1:0] ram_w32_l512_id4_1_rdata;
  wire [32-1:0] ram_w32_l512_id4_1_wdata;
  wire ram_w32_l512_id4_1_wenable;
  wire ram_w32_l512_id4_1_enable;
  assign ram_w32_l512_id4_0_wdata = 'hx;
  assign ram_w32_l512_id4_0_wenable = 0;

  ram_w32_l512_id4
  inst_ram_w32_l512_id4
  (
    .CLK(CLK),
    .ram_w32_l512_id4_0_addr(ram_w32_l512_id4_0_addr),
    .ram_w32_l512_id4_0_rdata(ram_w32_l512_id4_0_rdata),
    .ram_w32_l512_id4_0_wdata(ram_w32_l512_id4_0_wdata),
    .ram_w32_l512_id4_0_wenable(ram_w32_l512_id4_0_wenable),
    .ram_w32_l512_id4_0_enable(ram_w32_l512_id4_0_enable),
    .ram_w32_l512_id4_1_addr(ram_w32_l512_id4_1_addr),
    .ram_w32_l512_id4_1_rdata(ram_w32_l512_id4_1_rdata),
    .ram_w32_l512_id4_1_wdata(ram_w32_l512_id4_1_wdata),
    .ram_w32_l512_id4_1_wenable(ram_w32_l512_id4_1_wenable),
    .ram_w32_l512_id4_1_enable(ram_w32_l512_id4_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id5_0_addr;
  wire [32-1:0] ram_w32_l512_id5_0_rdata;
  wire [32-1:0] ram_w32_l512_id5_0_wdata;
  wire ram_w32_l512_id5_0_wenable;
  wire ram_w32_l512_id5_0_enable;
  wire [9-1:0] ram_w32_l512_id5_1_addr;
  wire [32-1:0] ram_w32_l512_id5_1_rdata;
  wire [32-1:0] ram_w32_l512_id5_1_wdata;
  wire ram_w32_l512_id5_1_wenable;
  wire ram_w32_l512_id5_1_enable;
  assign ram_w32_l512_id5_0_wdata = 'hx;
  assign ram_w32_l512_id5_0_wenable = 0;

  ram_w32_l512_id5
  inst_ram_w32_l512_id5
  (
    .CLK(CLK),
    .ram_w32_l512_id5_0_addr(ram_w32_l512_id5_0_addr),
    .ram_w32_l512_id5_0_rdata(ram_w32_l512_id5_0_rdata),
    .ram_w32_l512_id5_0_wdata(ram_w32_l512_id5_0_wdata),
    .ram_w32_l512_id5_0_wenable(ram_w32_l512_id5_0_wenable),
    .ram_w32_l512_id5_0_enable(ram_w32_l512_id5_0_enable),
    .ram_w32_l512_id5_1_addr(ram_w32_l512_id5_1_addr),
    .ram_w32_l512_id5_1_rdata(ram_w32_l512_id5_1_rdata),
    .ram_w32_l512_id5_1_wdata(ram_w32_l512_id5_1_wdata),
    .ram_w32_l512_id5_1_wenable(ram_w32_l512_id5_1_wenable),
    .ram_w32_l512_id5_1_enable(ram_w32_l512_id5_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id6_0_addr;
  wire [32-1:0] ram_w32_l512_id6_0_rdata;
  wire [32-1:0] ram_w32_l512_id6_0_wdata;
  wire ram_w32_l512_id6_0_wenable;
  wire ram_w32_l512_id6_0_enable;
  wire [9-1:0] ram_w32_l512_id6_1_addr;
  wire [32-1:0] ram_w32_l512_id6_1_rdata;
  wire [32-1:0] ram_w32_l512_id6_1_wdata;
  wire ram_w32_l512_id6_1_wenable;
  wire ram_w32_l512_id6_1_enable;
  assign ram_w32_l512_id6_0_wdata = 'hx;
  assign ram_w32_l512_id6_0_wenable = 0;

  ram_w32_l512_id6
  inst_ram_w32_l512_id6
  (
    .CLK(CLK),
    .ram_w32_l512_id6_0_addr(ram_w32_l512_id6_0_addr),
    .ram_w32_l512_id6_0_rdata(ram_w32_l512_id6_0_rdata),
    .ram_w32_l512_id6_0_wdata(ram_w32_l512_id6_0_wdata),
    .ram_w32_l512_id6_0_wenable(ram_w32_l512_id6_0_wenable),
    .ram_w32_l512_id6_0_enable(ram_w32_l512_id6_0_enable),
    .ram_w32_l512_id6_1_addr(ram_w32_l512_id6_1_addr),
    .ram_w32_l512_id6_1_rdata(ram_w32_l512_id6_1_rdata),
    .ram_w32_l512_id6_1_wdata(ram_w32_l512_id6_1_wdata),
    .ram_w32_l512_id6_1_wenable(ram_w32_l512_id6_1_wenable),
    .ram_w32_l512_id6_1_enable(ram_w32_l512_id6_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id7_0_addr;
  wire [32-1:0] ram_w32_l512_id7_0_rdata;
  wire [32-1:0] ram_w32_l512_id7_0_wdata;
  wire ram_w32_l512_id7_0_wenable;
  wire ram_w32_l512_id7_0_enable;
  wire [9-1:0] ram_w32_l512_id7_1_addr;
  wire [32-1:0] ram_w32_l512_id7_1_rdata;
  wire [32-1:0] ram_w32_l512_id7_1_wdata;
  wire ram_w32_l512_id7_1_wenable;
  wire ram_w32_l512_id7_1_enable;
  assign ram_w32_l512_id7_0_wdata = 'hx;
  assign ram_w32_l512_id7_0_wenable = 0;

  ram_w32_l512_id7
  inst_ram_w32_l512_id7
  (
    .CLK(CLK),
    .ram_w32_l512_id7_0_addr(ram_w32_l512_id7_0_addr),
    .ram_w32_l512_id7_0_rdata(ram_w32_l512_id7_0_rdata),
    .ram_w32_l512_id7_0_wdata(ram_w32_l512_id7_0_wdata),
    .ram_w32_l512_id7_0_wenable(ram_w32_l512_id7_0_wenable),
    .ram_w32_l512_id7_0_enable(ram_w32_l512_id7_0_enable),
    .ram_w32_l512_id7_1_addr(ram_w32_l512_id7_1_addr),
    .ram_w32_l512_id7_1_rdata(ram_w32_l512_id7_1_rdata),
    .ram_w32_l512_id7_1_wdata(ram_w32_l512_id7_1_wdata),
    .ram_w32_l512_id7_1_wenable(ram_w32_l512_id7_1_wenable),
    .ram_w32_l512_id7_1_enable(ram_w32_l512_id7_1_enable)
  );

  wire [9-1:0] ram_w32_l512_id8_0_addr;
  wire [32-1:0] ram_w32_l512_id8_0_rdata;
  wire [32-1:0] ram_w32_l512_id8_0_wdata;
  wire ram_w32_l512_id8_0_wenable;
  wire ram_w32_l512_id8_0_enable;
  wire [9-1:0] ram_w32_l512_id8_1_addr;
  wire [32-1:0] ram_w32_l512_id8_1_rdata;
  wire [32-1:0] ram_w32_l512_id8_1_wdata;
  wire ram_w32_l512_id8_1_wenable;
  wire ram_w32_l512_id8_1_enable;
  assign ram_w32_l512_id8_0_wdata = 'hx;
  assign ram_w32_l512_id8_0_wenable = 0;

  ram_w32_l512_id8
  inst_ram_w32_l512_id8
  (
    .CLK(CLK),
    .ram_w32_l512_id8_0_addr(ram_w32_l512_id8_0_addr),
    .ram_w32_l512_id8_0_rdata(ram_w32_l512_id8_0_rdata),
    .ram_w32_l512_id8_0_wdata(ram_w32_l512_id8_0_wdata),
    .ram_w32_l512_id8_0_wenable(ram_w32_l512_id8_0_wenable),
    .ram_w32_l512_id8_0_enable(ram_w32_l512_id8_0_enable),
    .ram_w32_l512_id8_1_addr(ram_w32_l512_id8_1_addr),
    .ram_w32_l512_id8_1_rdata(ram_w32_l512_id8_1_rdata),
    .ram_w32_l512_id8_1_wdata(ram_w32_l512_id8_1_wdata),
    .ram_w32_l512_id8_1_wenable(ram_w32_l512_id8_1_wenable),
    .ram_w32_l512_id8_1_enable(ram_w32_l512_id8_1_enable)
  );

  wire [8-1:0] ram_w32_l256_id0_0_addr;
  wire [32-1:0] ram_w32_l256_id0_0_rdata;
  wire [32-1:0] ram_w32_l256_id0_0_wdata;
  wire ram_w32_l256_id0_0_wenable;
  wire ram_w32_l256_id0_0_enable;
  wire [8-1:0] ram_w32_l256_id0_1_addr;
  wire [32-1:0] ram_w32_l256_id0_1_rdata;
  wire [32-1:0] ram_w32_l256_id0_1_wdata;
  wire ram_w32_l256_id0_1_wenable;
  wire ram_w32_l256_id0_1_enable;
  assign ram_w32_l256_id0_0_wdata = 'hx;
  assign ram_w32_l256_id0_0_wenable = 0;

  ram_w32_l256_id0
  inst_ram_w32_l256_id0
  (
    .CLK(CLK),
    .ram_w32_l256_id0_0_addr(ram_w32_l256_id0_0_addr),
    .ram_w32_l256_id0_0_rdata(ram_w32_l256_id0_0_rdata),
    .ram_w32_l256_id0_0_wdata(ram_w32_l256_id0_0_wdata),
    .ram_w32_l256_id0_0_wenable(ram_w32_l256_id0_0_wenable),
    .ram_w32_l256_id0_0_enable(ram_w32_l256_id0_0_enable),
    .ram_w32_l256_id0_1_addr(ram_w32_l256_id0_1_addr),
    .ram_w32_l256_id0_1_rdata(ram_w32_l256_id0_1_rdata),
    .ram_w32_l256_id0_1_wdata(ram_w32_l256_id0_1_wdata),
    .ram_w32_l256_id0_1_wenable(ram_w32_l256_id0_1_wenable),
    .ram_w32_l256_id0_1_enable(ram_w32_l256_id0_1_enable)
  );

  wire [8-1:0] ram_w32_l256_id1_0_addr;
  wire [32-1:0] ram_w32_l256_id1_0_rdata;
  wire [32-1:0] ram_w32_l256_id1_0_wdata;
  wire ram_w32_l256_id1_0_wenable;
  wire ram_w32_l256_id1_0_enable;
  wire [8-1:0] ram_w32_l256_id1_1_addr;
  wire [32-1:0] ram_w32_l256_id1_1_rdata;
  wire [32-1:0] ram_w32_l256_id1_1_wdata;
  wire ram_w32_l256_id1_1_wenable;
  wire ram_w32_l256_id1_1_enable;
  assign ram_w32_l256_id1_0_wdata = 'hx;
  assign ram_w32_l256_id1_0_wenable = 0;

  ram_w32_l256_id1
  inst_ram_w32_l256_id1
  (
    .CLK(CLK),
    .ram_w32_l256_id1_0_addr(ram_w32_l256_id1_0_addr),
    .ram_w32_l256_id1_0_rdata(ram_w32_l256_id1_0_rdata),
    .ram_w32_l256_id1_0_wdata(ram_w32_l256_id1_0_wdata),
    .ram_w32_l256_id1_0_wenable(ram_w32_l256_id1_0_wenable),
    .ram_w32_l256_id1_0_enable(ram_w32_l256_id1_0_enable),
    .ram_w32_l256_id1_1_addr(ram_w32_l256_id1_1_addr),
    .ram_w32_l256_id1_1_rdata(ram_w32_l256_id1_1_rdata),
    .ram_w32_l256_id1_1_wdata(ram_w32_l256_id1_1_wdata),
    .ram_w32_l256_id1_1_wenable(ram_w32_l256_id1_1_wenable),
    .ram_w32_l256_id1_1_enable(ram_w32_l256_id1_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id0_0_addr;
  wire [32-1:0] ram_w32_l128_id0_0_rdata;
  wire [32-1:0] ram_w32_l128_id0_0_wdata;
  wire ram_w32_l128_id0_0_wenable;
  wire ram_w32_l128_id0_0_enable;
  wire [7-1:0] ram_w32_l128_id0_1_addr;
  wire [32-1:0] ram_w32_l128_id0_1_rdata;
  wire [32-1:0] ram_w32_l128_id0_1_wdata;
  wire ram_w32_l128_id0_1_wenable;
  wire ram_w32_l128_id0_1_enable;

  ram_w32_l128_id0
  inst_ram_w32_l128_id0
  (
    .CLK(CLK),
    .ram_w32_l128_id0_0_addr(ram_w32_l128_id0_0_addr),
    .ram_w32_l128_id0_0_rdata(ram_w32_l128_id0_0_rdata),
    .ram_w32_l128_id0_0_wdata(ram_w32_l128_id0_0_wdata),
    .ram_w32_l128_id0_0_wenable(ram_w32_l128_id0_0_wenable),
    .ram_w32_l128_id0_0_enable(ram_w32_l128_id0_0_enable),
    .ram_w32_l128_id0_1_addr(ram_w32_l128_id0_1_addr),
    .ram_w32_l128_id0_1_rdata(ram_w32_l128_id0_1_rdata),
    .ram_w32_l128_id0_1_wdata(ram_w32_l128_id0_1_wdata),
    .ram_w32_l128_id0_1_wenable(ram_w32_l128_id0_1_wenable),
    .ram_w32_l128_id0_1_enable(ram_w32_l128_id0_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id1_0_addr;
  wire [32-1:0] ram_w32_l128_id1_0_rdata;
  wire [32-1:0] ram_w32_l128_id1_0_wdata;
  wire ram_w32_l128_id1_0_wenable;
  wire ram_w32_l128_id1_0_enable;
  wire [7-1:0] ram_w32_l128_id1_1_addr;
  wire [32-1:0] ram_w32_l128_id1_1_rdata;
  wire [32-1:0] ram_w32_l128_id1_1_wdata;
  wire ram_w32_l128_id1_1_wenable;
  wire ram_w32_l128_id1_1_enable;
  assign ram_w32_l128_id1_0_wdata = 'hx;
  assign ram_w32_l128_id1_0_wenable = 0;

  ram_w32_l128_id1
  inst_ram_w32_l128_id1
  (
    .CLK(CLK),
    .ram_w32_l128_id1_0_addr(ram_w32_l128_id1_0_addr),
    .ram_w32_l128_id1_0_rdata(ram_w32_l128_id1_0_rdata),
    .ram_w32_l128_id1_0_wdata(ram_w32_l128_id1_0_wdata),
    .ram_w32_l128_id1_0_wenable(ram_w32_l128_id1_0_wenable),
    .ram_w32_l128_id1_0_enable(ram_w32_l128_id1_0_enable),
    .ram_w32_l128_id1_1_addr(ram_w32_l128_id1_1_addr),
    .ram_w32_l128_id1_1_rdata(ram_w32_l128_id1_1_rdata),
    .ram_w32_l128_id1_1_wdata(ram_w32_l128_id1_1_wdata),
    .ram_w32_l128_id1_1_wenable(ram_w32_l128_id1_1_wenable),
    .ram_w32_l128_id1_1_enable(ram_w32_l128_id1_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id2_0_addr;
  wire [32-1:0] ram_w32_l128_id2_0_rdata;
  wire [32-1:0] ram_w32_l128_id2_0_wdata;
  wire ram_w32_l128_id2_0_wenable;
  wire ram_w32_l128_id2_0_enable;
  wire [7-1:0] ram_w32_l128_id2_1_addr;
  wire [32-1:0] ram_w32_l128_id2_1_rdata;
  wire [32-1:0] ram_w32_l128_id2_1_wdata;
  wire ram_w32_l128_id2_1_wenable;
  wire ram_w32_l128_id2_1_enable;
  assign ram_w32_l128_id2_0_wdata = 'hx;
  assign ram_w32_l128_id2_0_wenable = 0;

  ram_w32_l128_id2
  inst_ram_w32_l128_id2
  (
    .CLK(CLK),
    .ram_w32_l128_id2_0_addr(ram_w32_l128_id2_0_addr),
    .ram_w32_l128_id2_0_rdata(ram_w32_l128_id2_0_rdata),
    .ram_w32_l128_id2_0_wdata(ram_w32_l128_id2_0_wdata),
    .ram_w32_l128_id2_0_wenable(ram_w32_l128_id2_0_wenable),
    .ram_w32_l128_id2_0_enable(ram_w32_l128_id2_0_enable),
    .ram_w32_l128_id2_1_addr(ram_w32_l128_id2_1_addr),
    .ram_w32_l128_id2_1_rdata(ram_w32_l128_id2_1_rdata),
    .ram_w32_l128_id2_1_wdata(ram_w32_l128_id2_1_wdata),
    .ram_w32_l128_id2_1_wenable(ram_w32_l128_id2_1_wenable),
    .ram_w32_l128_id2_1_enable(ram_w32_l128_id2_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id3_0_addr;
  wire [32-1:0] ram_w32_l128_id3_0_rdata;
  wire [32-1:0] ram_w32_l128_id3_0_wdata;
  wire ram_w32_l128_id3_0_wenable;
  wire ram_w32_l128_id3_0_enable;
  wire [7-1:0] ram_w32_l128_id3_1_addr;
  wire [32-1:0] ram_w32_l128_id3_1_rdata;
  wire [32-1:0] ram_w32_l128_id3_1_wdata;
  wire ram_w32_l128_id3_1_wenable;
  wire ram_w32_l128_id3_1_enable;
  assign ram_w32_l128_id3_0_wdata = 'hx;
  assign ram_w32_l128_id3_0_wenable = 0;

  ram_w32_l128_id3
  inst_ram_w32_l128_id3
  (
    .CLK(CLK),
    .ram_w32_l128_id3_0_addr(ram_w32_l128_id3_0_addr),
    .ram_w32_l128_id3_0_rdata(ram_w32_l128_id3_0_rdata),
    .ram_w32_l128_id3_0_wdata(ram_w32_l128_id3_0_wdata),
    .ram_w32_l128_id3_0_wenable(ram_w32_l128_id3_0_wenable),
    .ram_w32_l128_id3_0_enable(ram_w32_l128_id3_0_enable),
    .ram_w32_l128_id3_1_addr(ram_w32_l128_id3_1_addr),
    .ram_w32_l128_id3_1_rdata(ram_w32_l128_id3_1_rdata),
    .ram_w32_l128_id3_1_wdata(ram_w32_l128_id3_1_wdata),
    .ram_w32_l128_id3_1_wenable(ram_w32_l128_id3_1_wenable),
    .ram_w32_l128_id3_1_enable(ram_w32_l128_id3_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id4_0_addr;
  wire [32-1:0] ram_w32_l128_id4_0_rdata;
  wire [32-1:0] ram_w32_l128_id4_0_wdata;
  wire ram_w32_l128_id4_0_wenable;
  wire ram_w32_l128_id4_0_enable;
  wire [7-1:0] ram_w32_l128_id4_1_addr;
  wire [32-1:0] ram_w32_l128_id4_1_rdata;
  wire [32-1:0] ram_w32_l128_id4_1_wdata;
  wire ram_w32_l128_id4_1_wenable;
  wire ram_w32_l128_id4_1_enable;
  assign ram_w32_l128_id4_0_wdata = 'hx;
  assign ram_w32_l128_id4_0_wenable = 0;

  ram_w32_l128_id4
  inst_ram_w32_l128_id4
  (
    .CLK(CLK),
    .ram_w32_l128_id4_0_addr(ram_w32_l128_id4_0_addr),
    .ram_w32_l128_id4_0_rdata(ram_w32_l128_id4_0_rdata),
    .ram_w32_l128_id4_0_wdata(ram_w32_l128_id4_0_wdata),
    .ram_w32_l128_id4_0_wenable(ram_w32_l128_id4_0_wenable),
    .ram_w32_l128_id4_0_enable(ram_w32_l128_id4_0_enable),
    .ram_w32_l128_id4_1_addr(ram_w32_l128_id4_1_addr),
    .ram_w32_l128_id4_1_rdata(ram_w32_l128_id4_1_rdata),
    .ram_w32_l128_id4_1_wdata(ram_w32_l128_id4_1_wdata),
    .ram_w32_l128_id4_1_wenable(ram_w32_l128_id4_1_wenable),
    .ram_w32_l128_id4_1_enable(ram_w32_l128_id4_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id5_0_addr;
  wire [32-1:0] ram_w32_l128_id5_0_rdata;
  wire [32-1:0] ram_w32_l128_id5_0_wdata;
  wire ram_w32_l128_id5_0_wenable;
  wire ram_w32_l128_id5_0_enable;
  wire [7-1:0] ram_w32_l128_id5_1_addr;
  wire [32-1:0] ram_w32_l128_id5_1_rdata;
  wire [32-1:0] ram_w32_l128_id5_1_wdata;
  wire ram_w32_l128_id5_1_wenable;
  wire ram_w32_l128_id5_1_enable;
  assign ram_w32_l128_id5_0_wdata = 'hx;
  assign ram_w32_l128_id5_0_wenable = 0;

  ram_w32_l128_id5
  inst_ram_w32_l128_id5
  (
    .CLK(CLK),
    .ram_w32_l128_id5_0_addr(ram_w32_l128_id5_0_addr),
    .ram_w32_l128_id5_0_rdata(ram_w32_l128_id5_0_rdata),
    .ram_w32_l128_id5_0_wdata(ram_w32_l128_id5_0_wdata),
    .ram_w32_l128_id5_0_wenable(ram_w32_l128_id5_0_wenable),
    .ram_w32_l128_id5_0_enable(ram_w32_l128_id5_0_enable),
    .ram_w32_l128_id5_1_addr(ram_w32_l128_id5_1_addr),
    .ram_w32_l128_id5_1_rdata(ram_w32_l128_id5_1_rdata),
    .ram_w32_l128_id5_1_wdata(ram_w32_l128_id5_1_wdata),
    .ram_w32_l128_id5_1_wenable(ram_w32_l128_id5_1_wenable),
    .ram_w32_l128_id5_1_enable(ram_w32_l128_id5_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id6_0_addr;
  wire [32-1:0] ram_w32_l128_id6_0_rdata;
  wire [32-1:0] ram_w32_l128_id6_0_wdata;
  wire ram_w32_l128_id6_0_wenable;
  wire ram_w32_l128_id6_0_enable;
  wire [7-1:0] ram_w32_l128_id6_1_addr;
  wire [32-1:0] ram_w32_l128_id6_1_rdata;
  wire [32-1:0] ram_w32_l128_id6_1_wdata;
  wire ram_w32_l128_id6_1_wenable;
  wire ram_w32_l128_id6_1_enable;
  assign ram_w32_l128_id6_0_wdata = 'hx;
  assign ram_w32_l128_id6_0_wenable = 0;

  ram_w32_l128_id6
  inst_ram_w32_l128_id6
  (
    .CLK(CLK),
    .ram_w32_l128_id6_0_addr(ram_w32_l128_id6_0_addr),
    .ram_w32_l128_id6_0_rdata(ram_w32_l128_id6_0_rdata),
    .ram_w32_l128_id6_0_wdata(ram_w32_l128_id6_0_wdata),
    .ram_w32_l128_id6_0_wenable(ram_w32_l128_id6_0_wenable),
    .ram_w32_l128_id6_0_enable(ram_w32_l128_id6_0_enable),
    .ram_w32_l128_id6_1_addr(ram_w32_l128_id6_1_addr),
    .ram_w32_l128_id6_1_rdata(ram_w32_l128_id6_1_rdata),
    .ram_w32_l128_id6_1_wdata(ram_w32_l128_id6_1_wdata),
    .ram_w32_l128_id6_1_wenable(ram_w32_l128_id6_1_wenable),
    .ram_w32_l128_id6_1_enable(ram_w32_l128_id6_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id7_0_addr;
  wire [32-1:0] ram_w32_l128_id7_0_rdata;
  wire [32-1:0] ram_w32_l128_id7_0_wdata;
  wire ram_w32_l128_id7_0_wenable;
  wire ram_w32_l128_id7_0_enable;
  wire [7-1:0] ram_w32_l128_id7_1_addr;
  wire [32-1:0] ram_w32_l128_id7_1_rdata;
  wire [32-1:0] ram_w32_l128_id7_1_wdata;
  wire ram_w32_l128_id7_1_wenable;
  wire ram_w32_l128_id7_1_enable;
  assign ram_w32_l128_id7_0_wdata = 'hx;
  assign ram_w32_l128_id7_0_wenable = 0;

  ram_w32_l128_id7
  inst_ram_w32_l128_id7
  (
    .CLK(CLK),
    .ram_w32_l128_id7_0_addr(ram_w32_l128_id7_0_addr),
    .ram_w32_l128_id7_0_rdata(ram_w32_l128_id7_0_rdata),
    .ram_w32_l128_id7_0_wdata(ram_w32_l128_id7_0_wdata),
    .ram_w32_l128_id7_0_wenable(ram_w32_l128_id7_0_wenable),
    .ram_w32_l128_id7_0_enable(ram_w32_l128_id7_0_enable),
    .ram_w32_l128_id7_1_addr(ram_w32_l128_id7_1_addr),
    .ram_w32_l128_id7_1_rdata(ram_w32_l128_id7_1_rdata),
    .ram_w32_l128_id7_1_wdata(ram_w32_l128_id7_1_wdata),
    .ram_w32_l128_id7_1_wenable(ram_w32_l128_id7_1_wenable),
    .ram_w32_l128_id7_1_enable(ram_w32_l128_id7_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id8_0_addr;
  wire [32-1:0] ram_w32_l128_id8_0_rdata;
  wire [32-1:0] ram_w32_l128_id8_0_wdata;
  wire ram_w32_l128_id8_0_wenable;
  wire ram_w32_l128_id8_0_enable;
  wire [7-1:0] ram_w32_l128_id8_1_addr;
  wire [32-1:0] ram_w32_l128_id8_1_rdata;
  wire [32-1:0] ram_w32_l128_id8_1_wdata;
  wire ram_w32_l128_id8_1_wenable;
  wire ram_w32_l128_id8_1_enable;
  assign ram_w32_l128_id8_0_wdata = 'hx;
  assign ram_w32_l128_id8_0_wenable = 0;

  ram_w32_l128_id8
  inst_ram_w32_l128_id8
  (
    .CLK(CLK),
    .ram_w32_l128_id8_0_addr(ram_w32_l128_id8_0_addr),
    .ram_w32_l128_id8_0_rdata(ram_w32_l128_id8_0_rdata),
    .ram_w32_l128_id8_0_wdata(ram_w32_l128_id8_0_wdata),
    .ram_w32_l128_id8_0_wenable(ram_w32_l128_id8_0_wenable),
    .ram_w32_l128_id8_0_enable(ram_w32_l128_id8_0_enable),
    .ram_w32_l128_id8_1_addr(ram_w32_l128_id8_1_addr),
    .ram_w32_l128_id8_1_rdata(ram_w32_l128_id8_1_rdata),
    .ram_w32_l128_id8_1_wdata(ram_w32_l128_id8_1_wdata),
    .ram_w32_l128_id8_1_wenable(ram_w32_l128_id8_1_wenable),
    .ram_w32_l128_id8_1_enable(ram_w32_l128_id8_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id9_0_addr;
  wire [32-1:0] ram_w32_l128_id9_0_rdata;
  wire [32-1:0] ram_w32_l128_id9_0_wdata;
  wire ram_w32_l128_id9_0_wenable;
  wire ram_w32_l128_id9_0_enable;
  wire [7-1:0] ram_w32_l128_id9_1_addr;
  wire [32-1:0] ram_w32_l128_id9_1_rdata;
  wire [32-1:0] ram_w32_l128_id9_1_wdata;
  wire ram_w32_l128_id9_1_wenable;
  wire ram_w32_l128_id9_1_enable;
  assign ram_w32_l128_id9_0_wdata = 'hx;
  assign ram_w32_l128_id9_0_wenable = 0;

  ram_w32_l128_id9
  inst_ram_w32_l128_id9
  (
    .CLK(CLK),
    .ram_w32_l128_id9_0_addr(ram_w32_l128_id9_0_addr),
    .ram_w32_l128_id9_0_rdata(ram_w32_l128_id9_0_rdata),
    .ram_w32_l128_id9_0_wdata(ram_w32_l128_id9_0_wdata),
    .ram_w32_l128_id9_0_wenable(ram_w32_l128_id9_0_wenable),
    .ram_w32_l128_id9_0_enable(ram_w32_l128_id9_0_enable),
    .ram_w32_l128_id9_1_addr(ram_w32_l128_id9_1_addr),
    .ram_w32_l128_id9_1_rdata(ram_w32_l128_id9_1_rdata),
    .ram_w32_l128_id9_1_wdata(ram_w32_l128_id9_1_wdata),
    .ram_w32_l128_id9_1_wenable(ram_w32_l128_id9_1_wenable),
    .ram_w32_l128_id9_1_enable(ram_w32_l128_id9_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id10_0_addr;
  wire [32-1:0] ram_w32_l128_id10_0_rdata;
  wire [32-1:0] ram_w32_l128_id10_0_wdata;
  wire ram_w32_l128_id10_0_wenable;
  wire ram_w32_l128_id10_0_enable;
  wire [7-1:0] ram_w32_l128_id10_1_addr;
  wire [32-1:0] ram_w32_l128_id10_1_rdata;
  wire [32-1:0] ram_w32_l128_id10_1_wdata;
  wire ram_w32_l128_id10_1_wenable;
  wire ram_w32_l128_id10_1_enable;
  assign ram_w32_l128_id10_0_wdata = 'hx;
  assign ram_w32_l128_id10_0_wenable = 0;

  ram_w32_l128_id10
  inst_ram_w32_l128_id10
  (
    .CLK(CLK),
    .ram_w32_l128_id10_0_addr(ram_w32_l128_id10_0_addr),
    .ram_w32_l128_id10_0_rdata(ram_w32_l128_id10_0_rdata),
    .ram_w32_l128_id10_0_wdata(ram_w32_l128_id10_0_wdata),
    .ram_w32_l128_id10_0_wenable(ram_w32_l128_id10_0_wenable),
    .ram_w32_l128_id10_0_enable(ram_w32_l128_id10_0_enable),
    .ram_w32_l128_id10_1_addr(ram_w32_l128_id10_1_addr),
    .ram_w32_l128_id10_1_rdata(ram_w32_l128_id10_1_rdata),
    .ram_w32_l128_id10_1_wdata(ram_w32_l128_id10_1_wdata),
    .ram_w32_l128_id10_1_wenable(ram_w32_l128_id10_1_wenable),
    .ram_w32_l128_id10_1_enable(ram_w32_l128_id10_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id11_0_addr;
  wire [32-1:0] ram_w32_l128_id11_0_rdata;
  wire [32-1:0] ram_w32_l128_id11_0_wdata;
  wire ram_w32_l128_id11_0_wenable;
  wire ram_w32_l128_id11_0_enable;
  wire [7-1:0] ram_w32_l128_id11_1_addr;
  wire [32-1:0] ram_w32_l128_id11_1_rdata;
  wire [32-1:0] ram_w32_l128_id11_1_wdata;
  wire ram_w32_l128_id11_1_wenable;
  wire ram_w32_l128_id11_1_enable;
  assign ram_w32_l128_id11_0_wdata = 'hx;
  assign ram_w32_l128_id11_0_wenable = 0;

  ram_w32_l128_id11
  inst_ram_w32_l128_id11
  (
    .CLK(CLK),
    .ram_w32_l128_id11_0_addr(ram_w32_l128_id11_0_addr),
    .ram_w32_l128_id11_0_rdata(ram_w32_l128_id11_0_rdata),
    .ram_w32_l128_id11_0_wdata(ram_w32_l128_id11_0_wdata),
    .ram_w32_l128_id11_0_wenable(ram_w32_l128_id11_0_wenable),
    .ram_w32_l128_id11_0_enable(ram_w32_l128_id11_0_enable),
    .ram_w32_l128_id11_1_addr(ram_w32_l128_id11_1_addr),
    .ram_w32_l128_id11_1_rdata(ram_w32_l128_id11_1_rdata),
    .ram_w32_l128_id11_1_wdata(ram_w32_l128_id11_1_wdata),
    .ram_w32_l128_id11_1_wenable(ram_w32_l128_id11_1_wenable),
    .ram_w32_l128_id11_1_enable(ram_w32_l128_id11_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id12_0_addr;
  wire [32-1:0] ram_w32_l128_id12_0_rdata;
  wire [32-1:0] ram_w32_l128_id12_0_wdata;
  wire ram_w32_l128_id12_0_wenable;
  wire ram_w32_l128_id12_0_enable;
  wire [7-1:0] ram_w32_l128_id12_1_addr;
  wire [32-1:0] ram_w32_l128_id12_1_rdata;
  wire [32-1:0] ram_w32_l128_id12_1_wdata;
  wire ram_w32_l128_id12_1_wenable;
  wire ram_w32_l128_id12_1_enable;
  assign ram_w32_l128_id12_0_wdata = 'hx;
  assign ram_w32_l128_id12_0_wenable = 0;

  ram_w32_l128_id12
  inst_ram_w32_l128_id12
  (
    .CLK(CLK),
    .ram_w32_l128_id12_0_addr(ram_w32_l128_id12_0_addr),
    .ram_w32_l128_id12_0_rdata(ram_w32_l128_id12_0_rdata),
    .ram_w32_l128_id12_0_wdata(ram_w32_l128_id12_0_wdata),
    .ram_w32_l128_id12_0_wenable(ram_w32_l128_id12_0_wenable),
    .ram_w32_l128_id12_0_enable(ram_w32_l128_id12_0_enable),
    .ram_w32_l128_id12_1_addr(ram_w32_l128_id12_1_addr),
    .ram_w32_l128_id12_1_rdata(ram_w32_l128_id12_1_rdata),
    .ram_w32_l128_id12_1_wdata(ram_w32_l128_id12_1_wdata),
    .ram_w32_l128_id12_1_wenable(ram_w32_l128_id12_1_wenable),
    .ram_w32_l128_id12_1_enable(ram_w32_l128_id12_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id13_0_addr;
  wire [32-1:0] ram_w32_l128_id13_0_rdata;
  wire [32-1:0] ram_w32_l128_id13_0_wdata;
  wire ram_w32_l128_id13_0_wenable;
  wire ram_w32_l128_id13_0_enable;
  wire [7-1:0] ram_w32_l128_id13_1_addr;
  wire [32-1:0] ram_w32_l128_id13_1_rdata;
  wire [32-1:0] ram_w32_l128_id13_1_wdata;
  wire ram_w32_l128_id13_1_wenable;
  wire ram_w32_l128_id13_1_enable;
  assign ram_w32_l128_id13_0_wdata = 'hx;
  assign ram_w32_l128_id13_0_wenable = 0;

  ram_w32_l128_id13
  inst_ram_w32_l128_id13
  (
    .CLK(CLK),
    .ram_w32_l128_id13_0_addr(ram_w32_l128_id13_0_addr),
    .ram_w32_l128_id13_0_rdata(ram_w32_l128_id13_0_rdata),
    .ram_w32_l128_id13_0_wdata(ram_w32_l128_id13_0_wdata),
    .ram_w32_l128_id13_0_wenable(ram_w32_l128_id13_0_wenable),
    .ram_w32_l128_id13_0_enable(ram_w32_l128_id13_0_enable),
    .ram_w32_l128_id13_1_addr(ram_w32_l128_id13_1_addr),
    .ram_w32_l128_id13_1_rdata(ram_w32_l128_id13_1_rdata),
    .ram_w32_l128_id13_1_wdata(ram_w32_l128_id13_1_wdata),
    .ram_w32_l128_id13_1_wenable(ram_w32_l128_id13_1_wenable),
    .ram_w32_l128_id13_1_enable(ram_w32_l128_id13_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id14_0_addr;
  wire [32-1:0] ram_w32_l128_id14_0_rdata;
  wire [32-1:0] ram_w32_l128_id14_0_wdata;
  wire ram_w32_l128_id14_0_wenable;
  wire ram_w32_l128_id14_0_enable;
  wire [7-1:0] ram_w32_l128_id14_1_addr;
  wire [32-1:0] ram_w32_l128_id14_1_rdata;
  wire [32-1:0] ram_w32_l128_id14_1_wdata;
  wire ram_w32_l128_id14_1_wenable;
  wire ram_w32_l128_id14_1_enable;
  assign ram_w32_l128_id14_0_wdata = 'hx;
  assign ram_w32_l128_id14_0_wenable = 0;

  ram_w32_l128_id14
  inst_ram_w32_l128_id14
  (
    .CLK(CLK),
    .ram_w32_l128_id14_0_addr(ram_w32_l128_id14_0_addr),
    .ram_w32_l128_id14_0_rdata(ram_w32_l128_id14_0_rdata),
    .ram_w32_l128_id14_0_wdata(ram_w32_l128_id14_0_wdata),
    .ram_w32_l128_id14_0_wenable(ram_w32_l128_id14_0_wenable),
    .ram_w32_l128_id14_0_enable(ram_w32_l128_id14_0_enable),
    .ram_w32_l128_id14_1_addr(ram_w32_l128_id14_1_addr),
    .ram_w32_l128_id14_1_rdata(ram_w32_l128_id14_1_rdata),
    .ram_w32_l128_id14_1_wdata(ram_w32_l128_id14_1_wdata),
    .ram_w32_l128_id14_1_wenable(ram_w32_l128_id14_1_wenable),
    .ram_w32_l128_id14_1_enable(ram_w32_l128_id14_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id15_0_addr;
  wire [32-1:0] ram_w32_l128_id15_0_rdata;
  wire [32-1:0] ram_w32_l128_id15_0_wdata;
  wire ram_w32_l128_id15_0_wenable;
  wire ram_w32_l128_id15_0_enable;
  wire [7-1:0] ram_w32_l128_id15_1_addr;
  wire [32-1:0] ram_w32_l128_id15_1_rdata;
  wire [32-1:0] ram_w32_l128_id15_1_wdata;
  wire ram_w32_l128_id15_1_wenable;
  wire ram_w32_l128_id15_1_enable;
  assign ram_w32_l128_id15_0_wdata = 'hx;
  assign ram_w32_l128_id15_0_wenable = 0;

  ram_w32_l128_id15
  inst_ram_w32_l128_id15
  (
    .CLK(CLK),
    .ram_w32_l128_id15_0_addr(ram_w32_l128_id15_0_addr),
    .ram_w32_l128_id15_0_rdata(ram_w32_l128_id15_0_rdata),
    .ram_w32_l128_id15_0_wdata(ram_w32_l128_id15_0_wdata),
    .ram_w32_l128_id15_0_wenable(ram_w32_l128_id15_0_wenable),
    .ram_w32_l128_id15_0_enable(ram_w32_l128_id15_0_enable),
    .ram_w32_l128_id15_1_addr(ram_w32_l128_id15_1_addr),
    .ram_w32_l128_id15_1_rdata(ram_w32_l128_id15_1_rdata),
    .ram_w32_l128_id15_1_wdata(ram_w32_l128_id15_1_wdata),
    .ram_w32_l128_id15_1_wenable(ram_w32_l128_id15_1_wenable),
    .ram_w32_l128_id15_1_enable(ram_w32_l128_id15_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id16_0_addr;
  wire [32-1:0] ram_w32_l128_id16_0_rdata;
  wire [32-1:0] ram_w32_l128_id16_0_wdata;
  wire ram_w32_l128_id16_0_wenable;
  wire ram_w32_l128_id16_0_enable;
  wire [7-1:0] ram_w32_l128_id16_1_addr;
  wire [32-1:0] ram_w32_l128_id16_1_rdata;
  wire [32-1:0] ram_w32_l128_id16_1_wdata;
  wire ram_w32_l128_id16_1_wenable;
  wire ram_w32_l128_id16_1_enable;
  assign ram_w32_l128_id16_0_wdata = 'hx;
  assign ram_w32_l128_id16_0_wenable = 0;

  ram_w32_l128_id16
  inst_ram_w32_l128_id16
  (
    .CLK(CLK),
    .ram_w32_l128_id16_0_addr(ram_w32_l128_id16_0_addr),
    .ram_w32_l128_id16_0_rdata(ram_w32_l128_id16_0_rdata),
    .ram_w32_l128_id16_0_wdata(ram_w32_l128_id16_0_wdata),
    .ram_w32_l128_id16_0_wenable(ram_w32_l128_id16_0_wenable),
    .ram_w32_l128_id16_0_enable(ram_w32_l128_id16_0_enable),
    .ram_w32_l128_id16_1_addr(ram_w32_l128_id16_1_addr),
    .ram_w32_l128_id16_1_rdata(ram_w32_l128_id16_1_rdata),
    .ram_w32_l128_id16_1_wdata(ram_w32_l128_id16_1_wdata),
    .ram_w32_l128_id16_1_wenable(ram_w32_l128_id16_1_wenable),
    .ram_w32_l128_id16_1_enable(ram_w32_l128_id16_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id17_0_addr;
  wire [32-1:0] ram_w32_l128_id17_0_rdata;
  wire [32-1:0] ram_w32_l128_id17_0_wdata;
  wire ram_w32_l128_id17_0_wenable;
  wire ram_w32_l128_id17_0_enable;
  wire [7-1:0] ram_w32_l128_id17_1_addr;
  wire [32-1:0] ram_w32_l128_id17_1_rdata;
  wire [32-1:0] ram_w32_l128_id17_1_wdata;
  wire ram_w32_l128_id17_1_wenable;
  wire ram_w32_l128_id17_1_enable;
  assign ram_w32_l128_id17_0_wdata = 'hx;
  assign ram_w32_l128_id17_0_wenable = 0;

  ram_w32_l128_id17
  inst_ram_w32_l128_id17
  (
    .CLK(CLK),
    .ram_w32_l128_id17_0_addr(ram_w32_l128_id17_0_addr),
    .ram_w32_l128_id17_0_rdata(ram_w32_l128_id17_0_rdata),
    .ram_w32_l128_id17_0_wdata(ram_w32_l128_id17_0_wdata),
    .ram_w32_l128_id17_0_wenable(ram_w32_l128_id17_0_wenable),
    .ram_w32_l128_id17_0_enable(ram_w32_l128_id17_0_enable),
    .ram_w32_l128_id17_1_addr(ram_w32_l128_id17_1_addr),
    .ram_w32_l128_id17_1_rdata(ram_w32_l128_id17_1_rdata),
    .ram_w32_l128_id17_1_wdata(ram_w32_l128_id17_1_wdata),
    .ram_w32_l128_id17_1_wenable(ram_w32_l128_id17_1_wenable),
    .ram_w32_l128_id17_1_enable(ram_w32_l128_id17_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id18_0_addr;
  wire [32-1:0] ram_w32_l128_id18_0_rdata;
  wire [32-1:0] ram_w32_l128_id18_0_wdata;
  wire ram_w32_l128_id18_0_wenable;
  wire ram_w32_l128_id18_0_enable;
  wire [7-1:0] ram_w32_l128_id18_1_addr;
  wire [32-1:0] ram_w32_l128_id18_1_rdata;
  wire [32-1:0] ram_w32_l128_id18_1_wdata;
  wire ram_w32_l128_id18_1_wenable;
  wire ram_w32_l128_id18_1_enable;
  assign ram_w32_l128_id18_0_wdata = 'hx;
  assign ram_w32_l128_id18_0_wenable = 0;

  ram_w32_l128_id18
  inst_ram_w32_l128_id18
  (
    .CLK(CLK),
    .ram_w32_l128_id18_0_addr(ram_w32_l128_id18_0_addr),
    .ram_w32_l128_id18_0_rdata(ram_w32_l128_id18_0_rdata),
    .ram_w32_l128_id18_0_wdata(ram_w32_l128_id18_0_wdata),
    .ram_w32_l128_id18_0_wenable(ram_w32_l128_id18_0_wenable),
    .ram_w32_l128_id18_0_enable(ram_w32_l128_id18_0_enable),
    .ram_w32_l128_id18_1_addr(ram_w32_l128_id18_1_addr),
    .ram_w32_l128_id18_1_rdata(ram_w32_l128_id18_1_rdata),
    .ram_w32_l128_id18_1_wdata(ram_w32_l128_id18_1_wdata),
    .ram_w32_l128_id18_1_wenable(ram_w32_l128_id18_1_wenable),
    .ram_w32_l128_id18_1_enable(ram_w32_l128_id18_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id19_0_addr;
  wire [32-1:0] ram_w32_l128_id19_0_rdata;
  wire [32-1:0] ram_w32_l128_id19_0_wdata;
  wire ram_w32_l128_id19_0_wenable;
  wire ram_w32_l128_id19_0_enable;
  wire [7-1:0] ram_w32_l128_id19_1_addr;
  wire [32-1:0] ram_w32_l128_id19_1_rdata;
  wire [32-1:0] ram_w32_l128_id19_1_wdata;
  wire ram_w32_l128_id19_1_wenable;
  wire ram_w32_l128_id19_1_enable;
  assign ram_w32_l128_id19_0_wdata = 'hx;
  assign ram_w32_l128_id19_0_wenable = 0;

  ram_w32_l128_id19
  inst_ram_w32_l128_id19
  (
    .CLK(CLK),
    .ram_w32_l128_id19_0_addr(ram_w32_l128_id19_0_addr),
    .ram_w32_l128_id19_0_rdata(ram_w32_l128_id19_0_rdata),
    .ram_w32_l128_id19_0_wdata(ram_w32_l128_id19_0_wdata),
    .ram_w32_l128_id19_0_wenable(ram_w32_l128_id19_0_wenable),
    .ram_w32_l128_id19_0_enable(ram_w32_l128_id19_0_enable),
    .ram_w32_l128_id19_1_addr(ram_w32_l128_id19_1_addr),
    .ram_w32_l128_id19_1_rdata(ram_w32_l128_id19_1_rdata),
    .ram_w32_l128_id19_1_wdata(ram_w32_l128_id19_1_wdata),
    .ram_w32_l128_id19_1_wenable(ram_w32_l128_id19_1_wenable),
    .ram_w32_l128_id19_1_enable(ram_w32_l128_id19_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id20_0_addr;
  wire [32-1:0] ram_w32_l128_id20_0_rdata;
  wire [32-1:0] ram_w32_l128_id20_0_wdata;
  wire ram_w32_l128_id20_0_wenable;
  wire ram_w32_l128_id20_0_enable;
  wire [7-1:0] ram_w32_l128_id20_1_addr;
  wire [32-1:0] ram_w32_l128_id20_1_rdata;
  wire [32-1:0] ram_w32_l128_id20_1_wdata;
  wire ram_w32_l128_id20_1_wenable;
  wire ram_w32_l128_id20_1_enable;
  assign ram_w32_l128_id20_1_wdata = 'hx;
  assign ram_w32_l128_id20_1_wenable = 0;

  ram_w32_l128_id20
  inst_ram_w32_l128_id20
  (
    .CLK(CLK),
    .ram_w32_l128_id20_0_addr(ram_w32_l128_id20_0_addr),
    .ram_w32_l128_id20_0_rdata(ram_w32_l128_id20_0_rdata),
    .ram_w32_l128_id20_0_wdata(ram_w32_l128_id20_0_wdata),
    .ram_w32_l128_id20_0_wenable(ram_w32_l128_id20_0_wenable),
    .ram_w32_l128_id20_0_enable(ram_w32_l128_id20_0_enable),
    .ram_w32_l128_id20_1_addr(ram_w32_l128_id20_1_addr),
    .ram_w32_l128_id20_1_rdata(ram_w32_l128_id20_1_rdata),
    .ram_w32_l128_id20_1_wdata(ram_w32_l128_id20_1_wdata),
    .ram_w32_l128_id20_1_wenable(ram_w32_l128_id20_1_wenable),
    .ram_w32_l128_id20_1_enable(ram_w32_l128_id20_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id21_0_addr;
  wire [32-1:0] ram_w32_l128_id21_0_rdata;
  wire [32-1:0] ram_w32_l128_id21_0_wdata;
  wire ram_w32_l128_id21_0_wenable;
  wire ram_w32_l128_id21_0_enable;
  wire [7-1:0] ram_w32_l128_id21_1_addr;
  wire [32-1:0] ram_w32_l128_id21_1_rdata;
  wire [32-1:0] ram_w32_l128_id21_1_wdata;
  wire ram_w32_l128_id21_1_wenable;
  wire ram_w32_l128_id21_1_enable;
  assign ram_w32_l128_id21_0_addr = 'hx;
  assign ram_w32_l128_id21_0_wdata = 'hx;
  assign ram_w32_l128_id21_0_wenable = 0;
  assign ram_w32_l128_id21_0_enable = 0;
  assign ram_w32_l128_id21_1_addr = 'hx;
  assign ram_w32_l128_id21_1_wdata = 'hx;
  assign ram_w32_l128_id21_1_wenable = 0;
  assign ram_w32_l128_id21_1_enable = 0;

  ram_w32_l128_id21
  inst_ram_w32_l128_id21
  (
    .CLK(CLK),
    .ram_w32_l128_id21_0_addr(ram_w32_l128_id21_0_addr),
    .ram_w32_l128_id21_0_rdata(ram_w32_l128_id21_0_rdata),
    .ram_w32_l128_id21_0_wdata(ram_w32_l128_id21_0_wdata),
    .ram_w32_l128_id21_0_wenable(ram_w32_l128_id21_0_wenable),
    .ram_w32_l128_id21_0_enable(ram_w32_l128_id21_0_enable),
    .ram_w32_l128_id21_1_addr(ram_w32_l128_id21_1_addr),
    .ram_w32_l128_id21_1_rdata(ram_w32_l128_id21_1_rdata),
    .ram_w32_l128_id21_1_wdata(ram_w32_l128_id21_1_wdata),
    .ram_w32_l128_id21_1_wenable(ram_w32_l128_id21_1_wenable),
    .ram_w32_l128_id21_1_enable(ram_w32_l128_id21_1_enable)
  );

  wire [6-1:0] cparam_conv2d_4_act_num_col;
  wire [6-1:0] cparam_conv2d_4_act_num_row;
  wire [7-1:0] cparam_conv2d_4_filter_num_och;
  wire [1-1:0] cparam_conv2d_4_bias_scala;
  wire [6-1:0] cparam_conv2d_4_bias_num;
  wire [1-1:0] cparam_conv2d_4_scale_scala;
  wire [6-1:0] cparam_conv2d_4_scale_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_mul_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_mul_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_sum_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_sum_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_out_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_out_num;
  wire [1-1:0] cparam_conv2d_4_cshamt_mul_value;
  wire [1-1:0] cparam_conv2d_4_cshamt_sum_value;
  wire [5-1:0] cparam_conv2d_4_cshamt_out_value;
  wire [1-1:0] cparam_conv2d_4_act_func_index;
  wire [6-1:0] cparam_conv2d_4_out_num_col;
  wire [6-1:0] cparam_conv2d_4_out_num_row;
  wire [1-1:0] cparam_conv2d_4_pad_col_left;
  wire [1-1:0] cparam_conv2d_4_pad_row_top;
  wire [5-1:0] cparam_conv2d_4_max_col_count;
  wire [5-1:0] cparam_conv2d_4_max_row_count;
  wire [1-1:0] cparam_conv2d_4_max_bat_count;
  wire [5-1:0] cparam_conv2d_4_max_och_count;
  wire [2-1:0] cparam_conv2d_4_och_count_step;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_0;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_1;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_2;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_0;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_1;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_2;
  wire [12-1:0] cparam_conv2d_4_act_row_step;
  wire [16-1:0] cparam_conv2d_4_act_bat_step;
  wire [10-1:0] cparam_conv2d_4_act_read_size;
  wire [6-1:0] cparam_conv2d_4_act_read_block;
  wire [8-1:0] cparam_conv2d_4_act_read_step;
  wire [13-1:0] cparam_conv2d_4_filter_base_step;
  wire [11-1:0] cparam_conv2d_4_filter_read_size;
  wire [6-1:0] cparam_conv2d_4_filter_read_block;
  wire [7-1:0] cparam_conv2d_4_filter_read_step;
  wire [1-1:0] cparam_conv2d_4_out_offset_values_0;
  wire [8-1:0] cparam_conv2d_4_out_col_step;
  wire [13-1:0] cparam_conv2d_4_out_row_step;
  wire [18-1:0] cparam_conv2d_4_out_bat_step;
  wire [4-1:0] cparam_conv2d_4_out_och_step;
  wire [2-1:0] cparam_conv2d_4_out_write_size;
  wire [2-1:0] cparam_conv2d_4_out_write_size_res;
  wire [1-1:0] cparam_conv2d_4_out_write_block;
  wire [1-1:0] cparam_conv2d_4_keep_filter;
  wire [1-1:0] cparam_conv2d_4_keep_input;
  wire [1-1:0] cparam_conv2d_4_data_stationary;
  wire [2-1:0] cparam_conv2d_4_stream_num_ops;
  wire [2-1:0] cparam_conv2d_4_stream_num_ops_res;
  wire [2-1:0] cparam_conv2d_4_stream_num_ops_par;
  wire [2-1:0] cparam_conv2d_4_stream_num_ops_res_par;
  wire [6-1:0] cparam_conv2d_4_stream_reduce_size;
  wire [6-1:0] cparam_conv2d_4_stream_aligned_reduce_size;
  wire [2-1:0] cparam_conv2d_4_stream_omit_mask;
  wire [2-1:0] cparam_conv2d_4_col_select_initval;
  wire [1-1:0] cparam_conv2d_4_stride_col_par_col;
  wire [1-1:0] cparam_conv2d_4_stride_row_par_row;
  wire [1-1:0] cparam_conv2d_4_stride_col_mod_filter_num;
  wire [2-1:0] cparam_conv2d_4_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_8;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_9;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_10;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_11;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_12;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_13;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_14;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_15;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_16;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_17;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_18;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_19;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_20;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_21;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_22;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_23;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_24;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_25;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_26;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_small;
  wire [6-1:0] cparam_conv2d_4_inc_act_laddr_large;
  wire [6-1:0] cparam_conv2d_4_inc_out_laddr_col;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_offset;
  wire signed [7-1:0] cparam_conv2d_4_stream_act_local_large_offset;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_2;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_1;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_2;
  wire [1-1:0] cparam_conv2d_4_inc_sync_out;
  wire [1-1:0] cparam_conv2d_4_inc_sync_out_res;
  reg [1-1:0] conv2d_4_control_param_index;
  assign cparam_conv2d_4_act_num_col = (conv2d_4_control_param_index == 0)? 32'h20 : 32'h10;
  assign cparam_conv2d_4_act_num_row = (conv2d_4_control_param_index == 0)? 32'h20 : 32'h10;
  assign cparam_conv2d_4_filter_num_och = (conv2d_4_control_param_index == 0)? 32'h40 : 32'h40;
  assign cparam_conv2d_4_bias_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_bias_num = (conv2d_4_control_param_index == 0)? 32'h20 : 32'h20;
  assign cparam_conv2d_4_scale_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_scale_num = (conv2d_4_control_param_index == 0)? 32'h20 : 32'h20;
  assign cparam_conv2d_4_vshamt_mul_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_mul_num = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_sum_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_sum_num = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_out_scala = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_vshamt_out_num = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_cshamt_mul_value = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_cshamt_sum_value = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_cshamt_out_value = (conv2d_4_control_param_index == 0)? 32'h11 : 32'h11;
  assign cparam_conv2d_4_act_func_index = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_out_num_col = (conv2d_4_control_param_index == 0)? 32'h20 : 32'h10;
  assign cparam_conv2d_4_out_num_row = (conv2d_4_control_param_index == 0)? 32'h20 : 32'h10;
  assign cparam_conv2d_4_pad_col_left = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_pad_row_top = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_max_col_count = (conv2d_4_control_param_index == 0)? 32'h1f : 32'hf;
  assign cparam_conv2d_4_max_row_count = (conv2d_4_control_param_index == 0)? 32'h1f : 32'hf;
  assign cparam_conv2d_4_max_bat_count = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_max_och_count = (conv2d_4_control_param_index == 0)? 32'h1e : 32'h1e;
  assign cparam_conv2d_4_och_count_step = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_dma_flag_conds_0 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_dma_flag_conds_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_dma_flag_conds_2 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_act_offset_values_0 = (conv2d_4_control_param_index == 0)? -32'sh100 : -32'sh800;
  assign cparam_conv2d_4_act_offset_values_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_act_offset_values_2 = (conv2d_4_control_param_index == 0)? 32'h100 : 32'h800;
  assign cparam_conv2d_4_act_row_step = (conv2d_4_control_param_index == 0)? 32'h100 : 32'h800;
  assign cparam_conv2d_4_act_bat_step = (conv2d_4_control_param_index == 0)? 32'h2000 : 32'h8000;
  assign cparam_conv2d_4_act_read_size = (conv2d_4_control_param_index == 0)? 32'h40 : 32'h200;
  assign cparam_conv2d_4_act_read_block = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h20;
  assign cparam_conv2d_4_act_read_step = (conv2d_4_control_param_index == 0)? 32'h16 : 32'hc0;
  assign cparam_conv2d_4_filter_base_step = (conv2d_4_control_param_index == 0)? 32'h120 : 32'h1200;
  assign cparam_conv2d_4_filter_read_size = (conv2d_4_control_param_index == 0)? 32'h48 : 32'h480;
  assign cparam_conv2d_4_filter_read_block = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h20;
  assign cparam_conv2d_4_filter_read_step = (conv2d_4_control_param_index == 0)? 32'h4 : 32'h40;
  assign cparam_conv2d_4_out_offset_values_0 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_out_col_step = (conv2d_4_control_param_index == 0)? 32'h80 : 32'h80;
  assign cparam_conv2d_4_out_row_step = (conv2d_4_control_param_index == 0)? 32'h1000 : 32'h800;
  assign cparam_conv2d_4_out_bat_step = (conv2d_4_control_param_index == 0)? 32'h20000 : 32'h8000;
  assign cparam_conv2d_4_out_och_step = (conv2d_4_control_param_index == 0)? 32'h8 : 32'h8;
  assign cparam_conv2d_4_out_write_size = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_out_write_size_res = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_out_write_block = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_keep_filter = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_keep_input = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h0;
  assign cparam_conv2d_4_data_stationary = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_num_ops = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_stream_num_ops_res = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_stream_num_ops_par = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_stream_num_ops_res_par = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_stream_reduce_size = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h20;
  assign cparam_conv2d_4_stream_aligned_reduce_size = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h20;
  assign cparam_conv2d_4_stream_omit_mask = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h0;
  assign cparam_conv2d_4_col_select_initval = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_stride_col_par_col = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_stride_row_par_row = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_stride_col_mod_filter_num = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_filter_num_col_minus_stride_col_mod = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h2;
  assign cparam_conv2d_4_inc_act_laddr_conds_0 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_2 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_3 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_4 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_5 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_6 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_7 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_8 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_9 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_10 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_11 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_12 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_13 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_14 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_15 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_16 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_17 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_18 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_19 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_20 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_21 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_22 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_conds_23 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_24 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_25 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_conds_26 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_act_laddr_small = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_inc_act_laddr_large = (conv2d_4_control_param_index == 0)? 32'h2 : 32'h20;
  assign cparam_conv2d_4_inc_out_laddr_col = (conv2d_4_control_param_index == 0)? 32'h20 : 32'h20;
  assign cparam_conv2d_4_stream_act_local_small_offset = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_large_offset = (conv2d_4_control_param_index == 0)? -32'sh2 : -32'sh20;
  assign cparam_conv2d_4_stream_act_local_small_flags_0 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_small_flags_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_small_flags_2 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_stream_act_local_large_flags_0 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_large_flags_1 = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_conv2d_4_stream_act_local_large_flags_2 = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_sync_out = (conv2d_4_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_conv2d_4_inc_sync_out_res = (conv2d_4_control_param_index == 0)? 32'h0 : 32'h0;
  wire [6-1:0] cparam_max_pool_serial_6_act_num_col;
  wire [6-1:0] cparam_max_pool_serial_6_act_num_row;
  wire [2-1:0] cparam_max_pool_serial_6_stride_col;
  wire [2-1:0] cparam_max_pool_serial_6_stride_row;
  wire [5-1:0] cparam_max_pool_serial_6_out_num_col;
  wire [5-1:0] cparam_max_pool_serial_6_out_num_row;
  wire [1-1:0] cparam_max_pool_serial_6_pad_col_left;
  wire [1-1:0] cparam_max_pool_serial_6_pad_row_top;
  wire [5-1:0] cparam_max_pool_serial_6_max_col_count;
  wire [5-1:0] cparam_max_pool_serial_6_max_row_count;
  wire [1-1:0] cparam_max_pool_serial_6_max_bat_count;
  wire signed [32-1:0] cparam_max_pool_serial_6_act_offset_values_0;
  wire signed [32-1:0] cparam_max_pool_serial_6_act_offset_values_1;
  wire [14-1:0] cparam_max_pool_serial_6_act_row_step;
  wire [18-1:0] cparam_max_pool_serial_6_act_bat_step;
  wire [11-1:0] cparam_max_pool_serial_6_act_read_size;
  wire [6-1:0] cparam_max_pool_serial_6_act_read_block;
  wire [12-1:0] cparam_max_pool_serial_6_out_row_step;
  wire [16-1:0] cparam_max_pool_serial_6_out_bat_step;
  wire [10-1:0] cparam_max_pool_serial_6_out_write_size;
  wire [6-1:0] cparam_max_pool_serial_6_stream_size;
  wire [1-1:0] cparam_max_pool_serial_6_col_select_initval;
  wire [1-1:0] cparam_max_pool_serial_6_stride_col_mod_ksize;
  wire [2-1:0] cparam_max_pool_serial_6_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_max_pool_serial_6_local_pad_offset;
  wire [7-1:0] cparam_max_pool_serial_6_inc_act_laddr;
  wire [6-1:0] cparam_max_pool_serial_6_inc_out_laddr;
  assign cparam_max_pool_serial_6_act_num_col = 32;
  assign cparam_max_pool_serial_6_act_num_row = 32;
  assign cparam_max_pool_serial_6_stride_col = 2;
  assign cparam_max_pool_serial_6_stride_row = 2;
  assign cparam_max_pool_serial_6_out_num_col = 16;
  assign cparam_max_pool_serial_6_out_num_row = 16;
  assign cparam_max_pool_serial_6_pad_col_left = 0;
  assign cparam_max_pool_serial_6_pad_row_top = 0;
  assign cparam_max_pool_serial_6_max_col_count = 29;
  assign cparam_max_pool_serial_6_max_row_count = 29;
  assign cparam_max_pool_serial_6_max_bat_count = 0;
  assign cparam_max_pool_serial_6_act_offset_values_0 = 0;
  assign cparam_max_pool_serial_6_act_offset_values_1 = 4096;
  assign cparam_max_pool_serial_6_act_row_step = 8192;
  assign cparam_max_pool_serial_6_act_bat_step = 131072;
  assign cparam_max_pool_serial_6_act_read_size = 1024;
  assign cparam_max_pool_serial_6_act_read_block = 32;
  assign cparam_max_pool_serial_6_out_row_step = 2048;
  assign cparam_max_pool_serial_6_out_bat_step = 32768;
  assign cparam_max_pool_serial_6_out_write_size = 512;
  assign cparam_max_pool_serial_6_stream_size = 32;
  assign cparam_max_pool_serial_6_col_select_initval = 0;
  assign cparam_max_pool_serial_6_stride_col_mod_ksize = 0;
  assign cparam_max_pool_serial_6_ksize_col_minus_stride_col_mod = 2;
  assign cparam_max_pool_serial_6_local_pad_offset = 0;
  assign cparam_max_pool_serial_6_inc_act_laddr = 64;
  assign cparam_max_pool_serial_6_inc_out_laddr = 32;
  wire [1-1:0] cparam_matmul_16_act_num_col;
  wire [1-1:0] cparam_matmul_16_act_num_row;
  wire [9-1:0] cparam_matmul_16_filter_num_och;
  wire [1-1:0] cparam_matmul_16_bias_scala;
  wire [8-1:0] cparam_matmul_16_bias_num;
  wire [1-1:0] cparam_matmul_16_scale_scala;
  wire [8-1:0] cparam_matmul_16_scale_num;
  wire [1-1:0] cparam_matmul_16_vshamt_mul_scala;
  wire [1-1:0] cparam_matmul_16_vshamt_mul_num;
  wire [1-1:0] cparam_matmul_16_vshamt_sum_scala;
  wire [1-1:0] cparam_matmul_16_vshamt_sum_num;
  wire [1-1:0] cparam_matmul_16_vshamt_out_scala;
  wire [1-1:0] cparam_matmul_16_vshamt_out_num;
  wire [1-1:0] cparam_matmul_16_cshamt_mul_value;
  wire [1-1:0] cparam_matmul_16_cshamt_sum_value;
  wire [5-1:0] cparam_matmul_16_cshamt_out_value;
  wire [1-1:0] cparam_matmul_16_act_func_index;
  wire [1-1:0] cparam_matmul_16_out_num_col;
  wire [1-1:0] cparam_matmul_16_out_num_row;
  wire [1-1:0] cparam_matmul_16_pad_col_left;
  wire [1-1:0] cparam_matmul_16_pad_row_top;
  wire [1-1:0] cparam_matmul_16_max_col_count;
  wire [1-1:0] cparam_matmul_16_max_row_count;
  wire [1-1:0] cparam_matmul_16_max_bat_count;
  wire [7-1:0] cparam_matmul_16_max_och_count;
  wire [7-1:0] cparam_matmul_16_och_count_step;
  wire [1-1:0] cparam_matmul_16_dma_flag_conds_0;
  wire signed [32-1:0] cparam_matmul_16_act_offset_values_0;
  wire [16-1:0] cparam_matmul_16_act_row_step;
  wire [16-1:0] cparam_matmul_16_act_bat_step;
  wire [14-1:0] cparam_matmul_16_act_read_size;
  wire [14-1:0] cparam_matmul_16_act_read_block;
  wire [14-1:0] cparam_matmul_16_act_read_step;
  wire [17-1:0] cparam_matmul_16_filter_base_step;
  wire [15-1:0] cparam_matmul_16_filter_read_size;
  wire [14-1:0] cparam_matmul_16_filter_read_block;
  wire [14-1:0] cparam_matmul_16_filter_read_step;
  wire [1-1:0] cparam_matmul_16_out_offset_values_0;
  wire [10-1:0] cparam_matmul_16_out_col_step;
  wire [10-1:0] cparam_matmul_16_out_row_step;
  wire [10-1:0] cparam_matmul_16_out_bat_step;
  wire [5-1:0] cparam_matmul_16_out_och_step;
  wire [3-1:0] cparam_matmul_16_out_write_size;
  wire [3-1:0] cparam_matmul_16_out_write_size_res;
  wire [3-1:0] cparam_matmul_16_out_write_block;
  wire [1-1:0] cparam_matmul_16_keep_filter;
  wire [1-1:0] cparam_matmul_16_keep_input;
  wire [1-1:0] cparam_matmul_16_data_stationary;
  wire [3-1:0] cparam_matmul_16_stream_num_ops;
  wire [3-1:0] cparam_matmul_16_stream_num_ops_res;
  wire [3-1:0] cparam_matmul_16_stream_num_ops_par;
  wire [3-1:0] cparam_matmul_16_stream_num_ops_res_par;
  wire [14-1:0] cparam_matmul_16_stream_reduce_size;
  wire [14-1:0] cparam_matmul_16_stream_aligned_reduce_size;
  wire [1-1:0] cparam_matmul_16_stream_omit_mask;
  wire [1-1:0] cparam_matmul_16_col_select_initval;
  wire [1-1:0] cparam_matmul_16_stride_col_par_col;
  wire [1-1:0] cparam_matmul_16_stride_row_par_row;
  wire [1-1:0] cparam_matmul_16_stride_col_mod_filter_num;
  wire [1-1:0] cparam_matmul_16_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_matmul_16_inc_act_laddr_conds_0;
  wire [14-1:0] cparam_matmul_16_inc_act_laddr_small;
  wire [14-1:0] cparam_matmul_16_inc_act_laddr_large;
  wire [8-1:0] cparam_matmul_16_inc_out_laddr_col;
  wire [1-1:0] cparam_matmul_16_stream_act_local_small_offset;
  wire [1-1:0] cparam_matmul_16_stream_act_local_large_offset;
  wire [1-1:0] cparam_matmul_16_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_matmul_16_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_matmul_16_inc_sync_out;
  wire [1-1:0] cparam_matmul_16_inc_sync_out_res;
  reg [1-1:0] matmul_16_control_param_index;
  assign cparam_matmul_16_act_num_col = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_act_num_row = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_filter_num_och = (matmul_16_control_param_index == 0)? 32'h100 : 32'ha;
  assign cparam_matmul_16_bias_scala = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_bias_num = (matmul_16_control_param_index == 0)? 32'h80 : 32'h5;
  assign cparam_matmul_16_scale_scala = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_scale_num = (matmul_16_control_param_index == 0)? 32'h80 : 32'h5;
  assign cparam_matmul_16_vshamt_mul_scala = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_vshamt_mul_num = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_vshamt_sum_scala = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_vshamt_sum_num = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_vshamt_out_scala = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_vshamt_out_num = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_cshamt_mul_value = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_cshamt_sum_value = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_cshamt_out_value = (matmul_16_control_param_index == 0)? 32'h11 : 32'h11;
  assign cparam_matmul_16_act_func_index = (matmul_16_control_param_index == 0)? 32'h0 : 32'h1;
  assign cparam_matmul_16_out_num_col = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_out_num_row = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_pad_col_left = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_pad_row_top = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_max_col_count = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_max_row_count = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_max_bat_count = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_max_och_count = (matmul_16_control_param_index == 0)? 32'h7f : 32'h0;
  assign cparam_matmul_16_och_count_step = (matmul_16_control_param_index == 0)? 32'h1 : 32'h40;
  assign cparam_matmul_16_dma_flag_conds_0 = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_act_offset_values_0 = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_act_row_step = (matmul_16_control_param_index == 0)? 32'h8000 : 32'h200;
  assign cparam_matmul_16_act_bat_step = (matmul_16_control_param_index == 0)? 32'h8000 : 32'h200;
  assign cparam_matmul_16_act_read_size = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_act_read_block = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_act_read_step = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_filter_base_step = (matmul_16_control_param_index == 0)? 32'h10000 : 32'h1400;
  assign cparam_matmul_16_filter_read_size = (matmul_16_control_param_index == 0)? 32'h4000 : 32'h500;
  assign cparam_matmul_16_filter_read_block = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_filter_read_step = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h280;
  assign cparam_matmul_16_out_offset_values_0 = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_out_col_step = (matmul_16_control_param_index == 0)? 32'h200 : 32'h14;
  assign cparam_matmul_16_out_row_step = (matmul_16_control_param_index == 0)? 32'h200 : 32'h14;
  assign cparam_matmul_16_out_bat_step = (matmul_16_control_param_index == 0)? 32'h200 : 32'h14;
  assign cparam_matmul_16_out_och_step = (matmul_16_control_param_index == 0)? 32'h4 : 32'h14;
  assign cparam_matmul_16_out_write_size = (matmul_16_control_param_index == 0)? 32'h1 : 32'h5;
  assign cparam_matmul_16_out_write_size_res = (matmul_16_control_param_index == 0)? 32'h1 : 32'h5;
  assign cparam_matmul_16_out_write_block = (matmul_16_control_param_index == 0)? 32'h0 : 32'h5;
  assign cparam_matmul_16_keep_filter = (matmul_16_control_param_index == 0)? 32'h0 : 32'h1;
  assign cparam_matmul_16_keep_input = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_data_stationary = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_stream_num_ops = (matmul_16_control_param_index == 0)? 32'h1 : 32'h5;
  assign cparam_matmul_16_stream_num_ops_res = (matmul_16_control_param_index == 0)? 32'h1 : 32'h5;
  assign cparam_matmul_16_stream_num_ops_par = (matmul_16_control_param_index == 0)? 32'h1 : 32'h5;
  assign cparam_matmul_16_stream_num_ops_res_par = (matmul_16_control_param_index == 0)? 32'h1 : 32'h5;
  assign cparam_matmul_16_stream_reduce_size = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_stream_aligned_reduce_size = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_stream_omit_mask = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_col_select_initval = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_stride_col_par_col = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_stride_row_par_row = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_stride_col_mod_filter_num = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_filter_num_col_minus_stride_col_mod = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_inc_act_laddr_conds_0 = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_inc_act_laddr_small = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_inc_act_laddr_large = (matmul_16_control_param_index == 0)? 32'h2000 : 32'h80;
  assign cparam_matmul_16_inc_out_laddr_col = (matmul_16_control_param_index == 0)? 32'h80 : 32'h5;
  assign cparam_matmul_16_stream_act_local_small_offset = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_stream_act_local_large_offset = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_stream_act_local_small_flags_0 = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_stream_act_local_large_flags_0 = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_16_inc_sync_out = (matmul_16_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_16_inc_sync_out_res = (matmul_16_control_param_index == 0)? 32'h0 : 32'h0;
  reg _acc_0_stream_ivalid;
  wire _acc_0_stream_oready;
  wire _acc_0_stream_internal_oready;
  assign _acc_0_stream_internal_oready = 1;
  reg [32-1:0] _acc_0_fsm;
  localparam _acc_0_fsm_init = 0;
  wire _acc_0_run_flag;
  assign _acc_0_run_flag = 0;
  reg _acc_0_source_start;
  wire _acc_0_source_stop;
  reg _acc_0_source_busy;
  wire _acc_0_sink_start;
  wire _acc_0_sink_stop;
  wire _acc_0_sink_busy;
  wire _acc_0_busy;
  reg _acc_0_busy_reg;
  wire _acc_0_is_root;
  reg _acc_0_x_idle;
  reg [33-1:0] _acc_0_x_source_count;
  reg [5-1:0] _acc_0_x_source_mode;
  reg [16-1:0] _acc_0_x_source_generator_id;
  reg [32-1:0] _acc_0_x_source_offset;
  reg [33-1:0] _acc_0_x_source_size;
  reg [32-1:0] _acc_0_x_source_stride;
  reg [32-1:0] _acc_0_x_source_offset_buf;
  reg [33-1:0] _acc_0_x_source_size_buf;
  reg [32-1:0] _acc_0_x_source_stride_buf;
  reg [8-1:0] _acc_0_x_source_sel;
  reg [32-1:0] _acc_0_x_source_ram_raddr;
  reg _acc_0_x_source_ram_renable;
  wire [64-1:0] _acc_0_x_source_ram_rdata;
  reg _acc_0_x_source_fifo_deq;
  wire [64-1:0] _acc_0_x_source_fifo_rdata;
  reg [64-1:0] _acc_0_x_source_empty_data;
  reg _acc_0_rshift_idle;
  reg [33-1:0] _acc_0_rshift_source_count;
  reg [5-1:0] _acc_0_rshift_source_mode;
  reg [16-1:0] _acc_0_rshift_source_generator_id;
  reg [32-1:0] _acc_0_rshift_source_offset;
  reg [33-1:0] _acc_0_rshift_source_size;
  reg [32-1:0] _acc_0_rshift_source_stride;
  reg [32-1:0] _acc_0_rshift_source_offset_buf;
  reg [33-1:0] _acc_0_rshift_source_size_buf;
  reg [32-1:0] _acc_0_rshift_source_stride_buf;
  reg [8-1:0] _acc_0_rshift_source_sel;
  reg [32-1:0] _acc_0_rshift_source_ram_raddr;
  reg _acc_0_rshift_source_ram_renable;
  wire [32-1:0] _acc_0_rshift_source_ram_rdata;
  reg _acc_0_rshift_source_fifo_deq;
  wire [32-1:0] _acc_0_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_0_rshift_source_empty_data;
  reg [32-1:0] _acc_0_size_next_parameter_data;
  reg [33-1:0] _acc_0_sum_sink_count;
  reg [5-1:0] _acc_0_sum_sink_mode;
  reg [16-1:0] _acc_0_sum_sink_generator_id;
  reg [32-1:0] _acc_0_sum_sink_offset;
  reg [33-1:0] _acc_0_sum_sink_size;
  reg [32-1:0] _acc_0_sum_sink_stride;
  reg [32-1:0] _acc_0_sum_sink_offset_buf;
  reg [33-1:0] _acc_0_sum_sink_size_buf;
  reg [32-1:0] _acc_0_sum_sink_stride_buf;
  reg [8-1:0] _acc_0_sum_sink_sel;
  reg [32-1:0] _acc_0_sum_sink_waddr;
  reg _acc_0_sum_sink_wenable;
  reg [64-1:0] _acc_0_sum_sink_wdata;
  reg _acc_0_sum_sink_fifo_enq;
  reg [64-1:0] _acc_0_sum_sink_fifo_wdata;
  reg [64-1:0] _acc_0_sum_sink_immediate;
  reg [33-1:0] _acc_0_valid_sink_count;
  reg [5-1:0] _acc_0_valid_sink_mode;
  reg [16-1:0] _acc_0_valid_sink_generator_id;
  reg [32-1:0] _acc_0_valid_sink_offset;
  reg [33-1:0] _acc_0_valid_sink_size;
  reg [32-1:0] _acc_0_valid_sink_stride;
  reg [32-1:0] _acc_0_valid_sink_offset_buf;
  reg [33-1:0] _acc_0_valid_sink_size_buf;
  reg [32-1:0] _acc_0_valid_sink_stride_buf;
  reg [8-1:0] _acc_0_valid_sink_sel;
  reg [32-1:0] _acc_0_valid_sink_waddr;
  reg _acc_0_valid_sink_wenable;
  reg [1-1:0] _acc_0_valid_sink_wdata;
  reg _acc_0_valid_sink_fifo_enq;
  reg [1-1:0] _acc_0_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_0_valid_sink_immediate;
  reg _acc_1_stream_ivalid;
  wire _acc_1_stream_oready;
  wire _acc_1_stream_internal_oready;
  assign _acc_1_stream_internal_oready = 1;
  reg [32-1:0] _acc_1_fsm;
  localparam _acc_1_fsm_init = 0;
  wire _acc_1_run_flag;
  assign _acc_1_run_flag = 0;
  reg _acc_1_source_start;
  wire _acc_1_source_stop;
  reg _acc_1_source_busy;
  wire _acc_1_sink_start;
  wire _acc_1_sink_stop;
  wire _acc_1_sink_busy;
  wire _acc_1_busy;
  reg _acc_1_busy_reg;
  wire _acc_1_is_root;
  reg _acc_1_x_idle;
  reg [33-1:0] _acc_1_x_source_count;
  reg [5-1:0] _acc_1_x_source_mode;
  reg [16-1:0] _acc_1_x_source_generator_id;
  reg [32-1:0] _acc_1_x_source_offset;
  reg [33-1:0] _acc_1_x_source_size;
  reg [32-1:0] _acc_1_x_source_stride;
  reg [32-1:0] _acc_1_x_source_offset_buf;
  reg [33-1:0] _acc_1_x_source_size_buf;
  reg [32-1:0] _acc_1_x_source_stride_buf;
  reg [8-1:0] _acc_1_x_source_sel;
  reg [32-1:0] _acc_1_x_source_ram_raddr;
  reg _acc_1_x_source_ram_renable;
  wire [64-1:0] _acc_1_x_source_ram_rdata;
  reg _acc_1_x_source_fifo_deq;
  wire [64-1:0] _acc_1_x_source_fifo_rdata;
  reg [64-1:0] _acc_1_x_source_empty_data;
  reg _acc_1_rshift_idle;
  reg [33-1:0] _acc_1_rshift_source_count;
  reg [5-1:0] _acc_1_rshift_source_mode;
  reg [16-1:0] _acc_1_rshift_source_generator_id;
  reg [32-1:0] _acc_1_rshift_source_offset;
  reg [33-1:0] _acc_1_rshift_source_size;
  reg [32-1:0] _acc_1_rshift_source_stride;
  reg [32-1:0] _acc_1_rshift_source_offset_buf;
  reg [33-1:0] _acc_1_rshift_source_size_buf;
  reg [32-1:0] _acc_1_rshift_source_stride_buf;
  reg [8-1:0] _acc_1_rshift_source_sel;
  reg [32-1:0] _acc_1_rshift_source_ram_raddr;
  reg _acc_1_rshift_source_ram_renable;
  wire [32-1:0] _acc_1_rshift_source_ram_rdata;
  reg _acc_1_rshift_source_fifo_deq;
  wire [32-1:0] _acc_1_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_1_rshift_source_empty_data;
  reg [32-1:0] _acc_1_size_next_parameter_data;
  reg [33-1:0] _acc_1_sum_sink_count;
  reg [5-1:0] _acc_1_sum_sink_mode;
  reg [16-1:0] _acc_1_sum_sink_generator_id;
  reg [32-1:0] _acc_1_sum_sink_offset;
  reg [33-1:0] _acc_1_sum_sink_size;
  reg [32-1:0] _acc_1_sum_sink_stride;
  reg [32-1:0] _acc_1_sum_sink_offset_buf;
  reg [33-1:0] _acc_1_sum_sink_size_buf;
  reg [32-1:0] _acc_1_sum_sink_stride_buf;
  reg [8-1:0] _acc_1_sum_sink_sel;
  reg [32-1:0] _acc_1_sum_sink_waddr;
  reg _acc_1_sum_sink_wenable;
  reg [64-1:0] _acc_1_sum_sink_wdata;
  reg _acc_1_sum_sink_fifo_enq;
  reg [64-1:0] _acc_1_sum_sink_fifo_wdata;
  reg [64-1:0] _acc_1_sum_sink_immediate;
  reg [33-1:0] _acc_1_valid_sink_count;
  reg [5-1:0] _acc_1_valid_sink_mode;
  reg [16-1:0] _acc_1_valid_sink_generator_id;
  reg [32-1:0] _acc_1_valid_sink_offset;
  reg [33-1:0] _acc_1_valid_sink_size;
  reg [32-1:0] _acc_1_valid_sink_stride;
  reg [32-1:0] _acc_1_valid_sink_offset_buf;
  reg [33-1:0] _acc_1_valid_sink_size_buf;
  reg [32-1:0] _acc_1_valid_sink_stride_buf;
  reg [8-1:0] _acc_1_valid_sink_sel;
  reg [32-1:0] _acc_1_valid_sink_waddr;
  reg _acc_1_valid_sink_wenable;
  reg [1-1:0] _acc_1_valid_sink_wdata;
  reg _acc_1_valid_sink_fifo_enq;
  reg [1-1:0] _acc_1_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_1_valid_sink_immediate;
  reg _add_tree_2_stream_ivalid;
  wire _add_tree_2_stream_oready;
  wire _add_tree_2_stream_internal_oready;
  assign _add_tree_2_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_2_fsm;
  localparam _add_tree_2_fsm_init = 0;
  wire _add_tree_2_run_flag;
  assign _add_tree_2_run_flag = 0;
  reg _add_tree_2_source_start;
  wire _add_tree_2_source_stop;
  reg _add_tree_2_source_busy;
  wire _add_tree_2_sink_start;
  wire _add_tree_2_sink_stop;
  wire _add_tree_2_sink_busy;
  wire _add_tree_2_busy;
  reg _add_tree_2_busy_reg;
  wire _add_tree_2_is_root;
  reg _add_tree_2_var0_idle;
  reg [33-1:0] _add_tree_2_var0_source_count;
  reg [5-1:0] _add_tree_2_var0_source_mode;
  reg [16-1:0] _add_tree_2_var0_source_generator_id;
  reg [32-1:0] _add_tree_2_var0_source_offset;
  reg [33-1:0] _add_tree_2_var0_source_size;
  reg [32-1:0] _add_tree_2_var0_source_stride;
  reg [32-1:0] _add_tree_2_var0_source_offset_buf;
  reg [33-1:0] _add_tree_2_var0_source_size_buf;
  reg [32-1:0] _add_tree_2_var0_source_stride_buf;
  reg [8-1:0] _add_tree_2_var0_source_sel;
  reg [32-1:0] _add_tree_2_var0_source_ram_raddr;
  reg _add_tree_2_var0_source_ram_renable;
  wire [64-1:0] _add_tree_2_var0_source_ram_rdata;
  reg _add_tree_2_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_2_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_2_var0_source_empty_data;
  reg _add_tree_2_var1_idle;
  reg [33-1:0] _add_tree_2_var1_source_count;
  reg [5-1:0] _add_tree_2_var1_source_mode;
  reg [16-1:0] _add_tree_2_var1_source_generator_id;
  reg [32-1:0] _add_tree_2_var1_source_offset;
  reg [33-1:0] _add_tree_2_var1_source_size;
  reg [32-1:0] _add_tree_2_var1_source_stride;
  reg [32-1:0] _add_tree_2_var1_source_offset_buf;
  reg [33-1:0] _add_tree_2_var1_source_size_buf;
  reg [32-1:0] _add_tree_2_var1_source_stride_buf;
  reg [8-1:0] _add_tree_2_var1_source_sel;
  reg [32-1:0] _add_tree_2_var1_source_ram_raddr;
  reg _add_tree_2_var1_source_ram_renable;
  wire [64-1:0] _add_tree_2_var1_source_ram_rdata;
  reg _add_tree_2_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_2_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_2_var1_source_empty_data;
  reg [33-1:0] _add_tree_2_sum_sink_count;
  reg [5-1:0] _add_tree_2_sum_sink_mode;
  reg [16-1:0] _add_tree_2_sum_sink_generator_id;
  reg [32-1:0] _add_tree_2_sum_sink_offset;
  reg [33-1:0] _add_tree_2_sum_sink_size;
  reg [32-1:0] _add_tree_2_sum_sink_stride;
  reg [32-1:0] _add_tree_2_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_2_sum_sink_size_buf;
  reg [32-1:0] _add_tree_2_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_2_sum_sink_sel;
  reg [32-1:0] _add_tree_2_sum_sink_waddr;
  reg _add_tree_2_sum_sink_wenable;
  reg [64-1:0] _add_tree_2_sum_sink_wdata;
  reg _add_tree_2_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_2_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_2_sum_sink_immediate;
  reg _add_tree_3_stream_ivalid;
  wire _add_tree_3_stream_oready;
  wire _add_tree_3_stream_internal_oready;
  assign _add_tree_3_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_3_fsm;
  localparam _add_tree_3_fsm_init = 0;
  wire _add_tree_3_run_flag;
  assign _add_tree_3_run_flag = 0;
  reg _add_tree_3_source_start;
  wire _add_tree_3_source_stop;
  reg _add_tree_3_source_busy;
  wire _add_tree_3_sink_start;
  wire _add_tree_3_sink_stop;
  wire _add_tree_3_sink_busy;
  wire _add_tree_3_busy;
  reg _add_tree_3_busy_reg;
  wire _add_tree_3_is_root;
  reg _add_tree_3_var0_idle;
  reg [33-1:0] _add_tree_3_var0_source_count;
  reg [5-1:0] _add_tree_3_var0_source_mode;
  reg [16-1:0] _add_tree_3_var0_source_generator_id;
  reg [32-1:0] _add_tree_3_var0_source_offset;
  reg [33-1:0] _add_tree_3_var0_source_size;
  reg [32-1:0] _add_tree_3_var0_source_stride;
  reg [32-1:0] _add_tree_3_var0_source_offset_buf;
  reg [33-1:0] _add_tree_3_var0_source_size_buf;
  reg [32-1:0] _add_tree_3_var0_source_stride_buf;
  reg [8-1:0] _add_tree_3_var0_source_sel;
  reg [32-1:0] _add_tree_3_var0_source_ram_raddr;
  reg _add_tree_3_var0_source_ram_renable;
  wire [64-1:0] _add_tree_3_var0_source_ram_rdata;
  reg _add_tree_3_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_3_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_3_var0_source_empty_data;
  reg _add_tree_3_var1_idle;
  reg [33-1:0] _add_tree_3_var1_source_count;
  reg [5-1:0] _add_tree_3_var1_source_mode;
  reg [16-1:0] _add_tree_3_var1_source_generator_id;
  reg [32-1:0] _add_tree_3_var1_source_offset;
  reg [33-1:0] _add_tree_3_var1_source_size;
  reg [32-1:0] _add_tree_3_var1_source_stride;
  reg [32-1:0] _add_tree_3_var1_source_offset_buf;
  reg [33-1:0] _add_tree_3_var1_source_size_buf;
  reg [32-1:0] _add_tree_3_var1_source_stride_buf;
  reg [8-1:0] _add_tree_3_var1_source_sel;
  reg [32-1:0] _add_tree_3_var1_source_ram_raddr;
  reg _add_tree_3_var1_source_ram_renable;
  wire [64-1:0] _add_tree_3_var1_source_ram_rdata;
  reg _add_tree_3_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_3_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_3_var1_source_empty_data;
  reg [33-1:0] _add_tree_3_sum_sink_count;
  reg [5-1:0] _add_tree_3_sum_sink_mode;
  reg [16-1:0] _add_tree_3_sum_sink_generator_id;
  reg [32-1:0] _add_tree_3_sum_sink_offset;
  reg [33-1:0] _add_tree_3_sum_sink_size;
  reg [32-1:0] _add_tree_3_sum_sink_stride;
  reg [32-1:0] _add_tree_3_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_3_sum_sink_size_buf;
  reg [32-1:0] _add_tree_3_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_3_sum_sink_sel;
  reg [32-1:0] _add_tree_3_sum_sink_waddr;
  reg _add_tree_3_sum_sink_wenable;
  reg [64-1:0] _add_tree_3_sum_sink_wdata;
  reg _add_tree_3_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_3_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_3_sum_sink_immediate;
  reg _add_tree_4_stream_ivalid;
  wire _add_tree_4_stream_oready;
  wire _add_tree_4_stream_internal_oready;
  assign _add_tree_4_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_4_fsm;
  localparam _add_tree_4_fsm_init = 0;
  wire _add_tree_4_run_flag;
  assign _add_tree_4_run_flag = 0;
  reg _add_tree_4_source_start;
  wire _add_tree_4_source_stop;
  reg _add_tree_4_source_busy;
  wire _add_tree_4_sink_start;
  wire _add_tree_4_sink_stop;
  wire _add_tree_4_sink_busy;
  wire _add_tree_4_busy;
  reg _add_tree_4_busy_reg;
  wire _add_tree_4_is_root;
  reg _add_tree_4_var0_idle;
  reg [33-1:0] _add_tree_4_var0_source_count;
  reg [5-1:0] _add_tree_4_var0_source_mode;
  reg [16-1:0] _add_tree_4_var0_source_generator_id;
  reg [32-1:0] _add_tree_4_var0_source_offset;
  reg [33-1:0] _add_tree_4_var0_source_size;
  reg [32-1:0] _add_tree_4_var0_source_stride;
  reg [32-1:0] _add_tree_4_var0_source_offset_buf;
  reg [33-1:0] _add_tree_4_var0_source_size_buf;
  reg [32-1:0] _add_tree_4_var0_source_stride_buf;
  reg [8-1:0] _add_tree_4_var0_source_sel;
  reg [32-1:0] _add_tree_4_var0_source_ram_raddr;
  reg _add_tree_4_var0_source_ram_renable;
  wire [64-1:0] _add_tree_4_var0_source_ram_rdata;
  reg _add_tree_4_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var0_source_empty_data;
  reg _add_tree_4_var1_idle;
  reg [33-1:0] _add_tree_4_var1_source_count;
  reg [5-1:0] _add_tree_4_var1_source_mode;
  reg [16-1:0] _add_tree_4_var1_source_generator_id;
  reg [32-1:0] _add_tree_4_var1_source_offset;
  reg [33-1:0] _add_tree_4_var1_source_size;
  reg [32-1:0] _add_tree_4_var1_source_stride;
  reg [32-1:0] _add_tree_4_var1_source_offset_buf;
  reg [33-1:0] _add_tree_4_var1_source_size_buf;
  reg [32-1:0] _add_tree_4_var1_source_stride_buf;
  reg [8-1:0] _add_tree_4_var1_source_sel;
  reg [32-1:0] _add_tree_4_var1_source_ram_raddr;
  reg _add_tree_4_var1_source_ram_renable;
  wire [64-1:0] _add_tree_4_var1_source_ram_rdata;
  reg _add_tree_4_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var1_source_empty_data;
  reg _add_tree_4_var2_idle;
  reg [33-1:0] _add_tree_4_var2_source_count;
  reg [5-1:0] _add_tree_4_var2_source_mode;
  reg [16-1:0] _add_tree_4_var2_source_generator_id;
  reg [32-1:0] _add_tree_4_var2_source_offset;
  reg [33-1:0] _add_tree_4_var2_source_size;
  reg [32-1:0] _add_tree_4_var2_source_stride;
  reg [32-1:0] _add_tree_4_var2_source_offset_buf;
  reg [33-1:0] _add_tree_4_var2_source_size_buf;
  reg [32-1:0] _add_tree_4_var2_source_stride_buf;
  reg [8-1:0] _add_tree_4_var2_source_sel;
  reg [32-1:0] _add_tree_4_var2_source_ram_raddr;
  reg _add_tree_4_var2_source_ram_renable;
  wire [64-1:0] _add_tree_4_var2_source_ram_rdata;
  reg _add_tree_4_var2_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var2_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var2_source_empty_data;
  reg _add_tree_4_var3_idle;
  reg [33-1:0] _add_tree_4_var3_source_count;
  reg [5-1:0] _add_tree_4_var3_source_mode;
  reg [16-1:0] _add_tree_4_var3_source_generator_id;
  reg [32-1:0] _add_tree_4_var3_source_offset;
  reg [33-1:0] _add_tree_4_var3_source_size;
  reg [32-1:0] _add_tree_4_var3_source_stride;
  reg [32-1:0] _add_tree_4_var3_source_offset_buf;
  reg [33-1:0] _add_tree_4_var3_source_size_buf;
  reg [32-1:0] _add_tree_4_var3_source_stride_buf;
  reg [8-1:0] _add_tree_4_var3_source_sel;
  reg [32-1:0] _add_tree_4_var3_source_ram_raddr;
  reg _add_tree_4_var3_source_ram_renable;
  wire [64-1:0] _add_tree_4_var3_source_ram_rdata;
  reg _add_tree_4_var3_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var3_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var3_source_empty_data;
  reg _add_tree_4_var4_idle;
  reg [33-1:0] _add_tree_4_var4_source_count;
  reg [5-1:0] _add_tree_4_var4_source_mode;
  reg [16-1:0] _add_tree_4_var4_source_generator_id;
  reg [32-1:0] _add_tree_4_var4_source_offset;
  reg [33-1:0] _add_tree_4_var4_source_size;
  reg [32-1:0] _add_tree_4_var4_source_stride;
  reg [32-1:0] _add_tree_4_var4_source_offset_buf;
  reg [33-1:0] _add_tree_4_var4_source_size_buf;
  reg [32-1:0] _add_tree_4_var4_source_stride_buf;
  reg [8-1:0] _add_tree_4_var4_source_sel;
  reg [32-1:0] _add_tree_4_var4_source_ram_raddr;
  reg _add_tree_4_var4_source_ram_renable;
  wire [64-1:0] _add_tree_4_var4_source_ram_rdata;
  reg _add_tree_4_var4_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var4_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var4_source_empty_data;
  reg _add_tree_4_var5_idle;
  reg [33-1:0] _add_tree_4_var5_source_count;
  reg [5-1:0] _add_tree_4_var5_source_mode;
  reg [16-1:0] _add_tree_4_var5_source_generator_id;
  reg [32-1:0] _add_tree_4_var5_source_offset;
  reg [33-1:0] _add_tree_4_var5_source_size;
  reg [32-1:0] _add_tree_4_var5_source_stride;
  reg [32-1:0] _add_tree_4_var5_source_offset_buf;
  reg [33-1:0] _add_tree_4_var5_source_size_buf;
  reg [32-1:0] _add_tree_4_var5_source_stride_buf;
  reg [8-1:0] _add_tree_4_var5_source_sel;
  reg [32-1:0] _add_tree_4_var5_source_ram_raddr;
  reg _add_tree_4_var5_source_ram_renable;
  wire [64-1:0] _add_tree_4_var5_source_ram_rdata;
  reg _add_tree_4_var5_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var5_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var5_source_empty_data;
  reg _add_tree_4_var6_idle;
  reg [33-1:0] _add_tree_4_var6_source_count;
  reg [5-1:0] _add_tree_4_var6_source_mode;
  reg [16-1:0] _add_tree_4_var6_source_generator_id;
  reg [32-1:0] _add_tree_4_var6_source_offset;
  reg [33-1:0] _add_tree_4_var6_source_size;
  reg [32-1:0] _add_tree_4_var6_source_stride;
  reg [32-1:0] _add_tree_4_var6_source_offset_buf;
  reg [33-1:0] _add_tree_4_var6_source_size_buf;
  reg [32-1:0] _add_tree_4_var6_source_stride_buf;
  reg [8-1:0] _add_tree_4_var6_source_sel;
  reg [32-1:0] _add_tree_4_var6_source_ram_raddr;
  reg _add_tree_4_var6_source_ram_renable;
  wire [64-1:0] _add_tree_4_var6_source_ram_rdata;
  reg _add_tree_4_var6_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var6_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var6_source_empty_data;
  reg _add_tree_4_var7_idle;
  reg [33-1:0] _add_tree_4_var7_source_count;
  reg [5-1:0] _add_tree_4_var7_source_mode;
  reg [16-1:0] _add_tree_4_var7_source_generator_id;
  reg [32-1:0] _add_tree_4_var7_source_offset;
  reg [33-1:0] _add_tree_4_var7_source_size;
  reg [32-1:0] _add_tree_4_var7_source_stride;
  reg [32-1:0] _add_tree_4_var7_source_offset_buf;
  reg [33-1:0] _add_tree_4_var7_source_size_buf;
  reg [32-1:0] _add_tree_4_var7_source_stride_buf;
  reg [8-1:0] _add_tree_4_var7_source_sel;
  reg [32-1:0] _add_tree_4_var7_source_ram_raddr;
  reg _add_tree_4_var7_source_ram_renable;
  wire [64-1:0] _add_tree_4_var7_source_ram_rdata;
  reg _add_tree_4_var7_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var7_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var7_source_empty_data;
  reg _add_tree_4_var8_idle;
  reg [33-1:0] _add_tree_4_var8_source_count;
  reg [5-1:0] _add_tree_4_var8_source_mode;
  reg [16-1:0] _add_tree_4_var8_source_generator_id;
  reg [32-1:0] _add_tree_4_var8_source_offset;
  reg [33-1:0] _add_tree_4_var8_source_size;
  reg [32-1:0] _add_tree_4_var8_source_stride;
  reg [32-1:0] _add_tree_4_var8_source_offset_buf;
  reg [33-1:0] _add_tree_4_var8_source_size_buf;
  reg [32-1:0] _add_tree_4_var8_source_stride_buf;
  reg [8-1:0] _add_tree_4_var8_source_sel;
  reg [32-1:0] _add_tree_4_var8_source_ram_raddr;
  reg _add_tree_4_var8_source_ram_renable;
  wire [64-1:0] _add_tree_4_var8_source_ram_rdata;
  reg _add_tree_4_var8_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var8_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var8_source_empty_data;
  reg _add_tree_4_var9_idle;
  reg [33-1:0] _add_tree_4_var9_source_count;
  reg [5-1:0] _add_tree_4_var9_source_mode;
  reg [16-1:0] _add_tree_4_var9_source_generator_id;
  reg [32-1:0] _add_tree_4_var9_source_offset;
  reg [33-1:0] _add_tree_4_var9_source_size;
  reg [32-1:0] _add_tree_4_var9_source_stride;
  reg [32-1:0] _add_tree_4_var9_source_offset_buf;
  reg [33-1:0] _add_tree_4_var9_source_size_buf;
  reg [32-1:0] _add_tree_4_var9_source_stride_buf;
  reg [8-1:0] _add_tree_4_var9_source_sel;
  reg [32-1:0] _add_tree_4_var9_source_ram_raddr;
  reg _add_tree_4_var9_source_ram_renable;
  wire [64-1:0] _add_tree_4_var9_source_ram_rdata;
  reg _add_tree_4_var9_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var9_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var9_source_empty_data;
  reg _add_tree_4_var10_idle;
  reg [33-1:0] _add_tree_4_var10_source_count;
  reg [5-1:0] _add_tree_4_var10_source_mode;
  reg [16-1:0] _add_tree_4_var10_source_generator_id;
  reg [32-1:0] _add_tree_4_var10_source_offset;
  reg [33-1:0] _add_tree_4_var10_source_size;
  reg [32-1:0] _add_tree_4_var10_source_stride;
  reg [32-1:0] _add_tree_4_var10_source_offset_buf;
  reg [33-1:0] _add_tree_4_var10_source_size_buf;
  reg [32-1:0] _add_tree_4_var10_source_stride_buf;
  reg [8-1:0] _add_tree_4_var10_source_sel;
  reg [32-1:0] _add_tree_4_var10_source_ram_raddr;
  reg _add_tree_4_var10_source_ram_renable;
  wire [64-1:0] _add_tree_4_var10_source_ram_rdata;
  reg _add_tree_4_var10_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var10_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var10_source_empty_data;
  reg _add_tree_4_var11_idle;
  reg [33-1:0] _add_tree_4_var11_source_count;
  reg [5-1:0] _add_tree_4_var11_source_mode;
  reg [16-1:0] _add_tree_4_var11_source_generator_id;
  reg [32-1:0] _add_tree_4_var11_source_offset;
  reg [33-1:0] _add_tree_4_var11_source_size;
  reg [32-1:0] _add_tree_4_var11_source_stride;
  reg [32-1:0] _add_tree_4_var11_source_offset_buf;
  reg [33-1:0] _add_tree_4_var11_source_size_buf;
  reg [32-1:0] _add_tree_4_var11_source_stride_buf;
  reg [8-1:0] _add_tree_4_var11_source_sel;
  reg [32-1:0] _add_tree_4_var11_source_ram_raddr;
  reg _add_tree_4_var11_source_ram_renable;
  wire [64-1:0] _add_tree_4_var11_source_ram_rdata;
  reg _add_tree_4_var11_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var11_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var11_source_empty_data;
  reg _add_tree_4_var12_idle;
  reg [33-1:0] _add_tree_4_var12_source_count;
  reg [5-1:0] _add_tree_4_var12_source_mode;
  reg [16-1:0] _add_tree_4_var12_source_generator_id;
  reg [32-1:0] _add_tree_4_var12_source_offset;
  reg [33-1:0] _add_tree_4_var12_source_size;
  reg [32-1:0] _add_tree_4_var12_source_stride;
  reg [32-1:0] _add_tree_4_var12_source_offset_buf;
  reg [33-1:0] _add_tree_4_var12_source_size_buf;
  reg [32-1:0] _add_tree_4_var12_source_stride_buf;
  reg [8-1:0] _add_tree_4_var12_source_sel;
  reg [32-1:0] _add_tree_4_var12_source_ram_raddr;
  reg _add_tree_4_var12_source_ram_renable;
  wire [64-1:0] _add_tree_4_var12_source_ram_rdata;
  reg _add_tree_4_var12_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var12_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var12_source_empty_data;
  reg _add_tree_4_var13_idle;
  reg [33-1:0] _add_tree_4_var13_source_count;
  reg [5-1:0] _add_tree_4_var13_source_mode;
  reg [16-1:0] _add_tree_4_var13_source_generator_id;
  reg [32-1:0] _add_tree_4_var13_source_offset;
  reg [33-1:0] _add_tree_4_var13_source_size;
  reg [32-1:0] _add_tree_4_var13_source_stride;
  reg [32-1:0] _add_tree_4_var13_source_offset_buf;
  reg [33-1:0] _add_tree_4_var13_source_size_buf;
  reg [32-1:0] _add_tree_4_var13_source_stride_buf;
  reg [8-1:0] _add_tree_4_var13_source_sel;
  reg [32-1:0] _add_tree_4_var13_source_ram_raddr;
  reg _add_tree_4_var13_source_ram_renable;
  wire [64-1:0] _add_tree_4_var13_source_ram_rdata;
  reg _add_tree_4_var13_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var13_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var13_source_empty_data;
  reg _add_tree_4_var14_idle;
  reg [33-1:0] _add_tree_4_var14_source_count;
  reg [5-1:0] _add_tree_4_var14_source_mode;
  reg [16-1:0] _add_tree_4_var14_source_generator_id;
  reg [32-1:0] _add_tree_4_var14_source_offset;
  reg [33-1:0] _add_tree_4_var14_source_size;
  reg [32-1:0] _add_tree_4_var14_source_stride;
  reg [32-1:0] _add_tree_4_var14_source_offset_buf;
  reg [33-1:0] _add_tree_4_var14_source_size_buf;
  reg [32-1:0] _add_tree_4_var14_source_stride_buf;
  reg [8-1:0] _add_tree_4_var14_source_sel;
  reg [32-1:0] _add_tree_4_var14_source_ram_raddr;
  reg _add_tree_4_var14_source_ram_renable;
  wire [64-1:0] _add_tree_4_var14_source_ram_rdata;
  reg _add_tree_4_var14_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var14_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var14_source_empty_data;
  reg _add_tree_4_var15_idle;
  reg [33-1:0] _add_tree_4_var15_source_count;
  reg [5-1:0] _add_tree_4_var15_source_mode;
  reg [16-1:0] _add_tree_4_var15_source_generator_id;
  reg [32-1:0] _add_tree_4_var15_source_offset;
  reg [33-1:0] _add_tree_4_var15_source_size;
  reg [32-1:0] _add_tree_4_var15_source_stride;
  reg [32-1:0] _add_tree_4_var15_source_offset_buf;
  reg [33-1:0] _add_tree_4_var15_source_size_buf;
  reg [32-1:0] _add_tree_4_var15_source_stride_buf;
  reg [8-1:0] _add_tree_4_var15_source_sel;
  reg [32-1:0] _add_tree_4_var15_source_ram_raddr;
  reg _add_tree_4_var15_source_ram_renable;
  wire [64-1:0] _add_tree_4_var15_source_ram_rdata;
  reg _add_tree_4_var15_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var15_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var15_source_empty_data;
  reg _add_tree_4_var16_idle;
  reg [33-1:0] _add_tree_4_var16_source_count;
  reg [5-1:0] _add_tree_4_var16_source_mode;
  reg [16-1:0] _add_tree_4_var16_source_generator_id;
  reg [32-1:0] _add_tree_4_var16_source_offset;
  reg [33-1:0] _add_tree_4_var16_source_size;
  reg [32-1:0] _add_tree_4_var16_source_stride;
  reg [32-1:0] _add_tree_4_var16_source_offset_buf;
  reg [33-1:0] _add_tree_4_var16_source_size_buf;
  reg [32-1:0] _add_tree_4_var16_source_stride_buf;
  reg [8-1:0] _add_tree_4_var16_source_sel;
  reg [32-1:0] _add_tree_4_var16_source_ram_raddr;
  reg _add_tree_4_var16_source_ram_renable;
  wire [64-1:0] _add_tree_4_var16_source_ram_rdata;
  reg _add_tree_4_var16_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var16_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var16_source_empty_data;
  reg _add_tree_4_var17_idle;
  reg [33-1:0] _add_tree_4_var17_source_count;
  reg [5-1:0] _add_tree_4_var17_source_mode;
  reg [16-1:0] _add_tree_4_var17_source_generator_id;
  reg [32-1:0] _add_tree_4_var17_source_offset;
  reg [33-1:0] _add_tree_4_var17_source_size;
  reg [32-1:0] _add_tree_4_var17_source_stride;
  reg [32-1:0] _add_tree_4_var17_source_offset_buf;
  reg [33-1:0] _add_tree_4_var17_source_size_buf;
  reg [32-1:0] _add_tree_4_var17_source_stride_buf;
  reg [8-1:0] _add_tree_4_var17_source_sel;
  reg [32-1:0] _add_tree_4_var17_source_ram_raddr;
  reg _add_tree_4_var17_source_ram_renable;
  wire [64-1:0] _add_tree_4_var17_source_ram_rdata;
  reg _add_tree_4_var17_source_fifo_deq;
  wire [64-1:0] _add_tree_4_var17_source_fifo_rdata;
  reg [64-1:0] _add_tree_4_var17_source_empty_data;
  reg [33-1:0] _add_tree_4_sum_sink_count;
  reg [5-1:0] _add_tree_4_sum_sink_mode;
  reg [16-1:0] _add_tree_4_sum_sink_generator_id;
  reg [32-1:0] _add_tree_4_sum_sink_offset;
  reg [33-1:0] _add_tree_4_sum_sink_size;
  reg [32-1:0] _add_tree_4_sum_sink_stride;
  reg [32-1:0] _add_tree_4_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_4_sum_sink_size_buf;
  reg [32-1:0] _add_tree_4_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_4_sum_sink_sel;
  reg [32-1:0] _add_tree_4_sum_sink_waddr;
  reg _add_tree_4_sum_sink_wenable;
  reg [64-1:0] _add_tree_4_sum_sink_wdata;
  reg _add_tree_4_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_4_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_4_sum_sink_immediate;
  reg _add_tree_5_stream_ivalid;
  wire _add_tree_5_stream_oready;
  wire _add_tree_5_stream_internal_oready;
  assign _add_tree_5_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_5_fsm;
  localparam _add_tree_5_fsm_init = 0;
  wire _add_tree_5_run_flag;
  assign _add_tree_5_run_flag = 0;
  reg _add_tree_5_source_start;
  wire _add_tree_5_source_stop;
  reg _add_tree_5_source_busy;
  wire _add_tree_5_sink_start;
  wire _add_tree_5_sink_stop;
  wire _add_tree_5_sink_busy;
  wire _add_tree_5_busy;
  reg _add_tree_5_busy_reg;
  wire _add_tree_5_is_root;
  reg _add_tree_5_var0_idle;
  reg [33-1:0] _add_tree_5_var0_source_count;
  reg [5-1:0] _add_tree_5_var0_source_mode;
  reg [16-1:0] _add_tree_5_var0_source_generator_id;
  reg [32-1:0] _add_tree_5_var0_source_offset;
  reg [33-1:0] _add_tree_5_var0_source_size;
  reg [32-1:0] _add_tree_5_var0_source_stride;
  reg [32-1:0] _add_tree_5_var0_source_offset_buf;
  reg [33-1:0] _add_tree_5_var0_source_size_buf;
  reg [32-1:0] _add_tree_5_var0_source_stride_buf;
  reg [8-1:0] _add_tree_5_var0_source_sel;
  reg [32-1:0] _add_tree_5_var0_source_ram_raddr;
  reg _add_tree_5_var0_source_ram_renable;
  wire [64-1:0] _add_tree_5_var0_source_ram_rdata;
  reg _add_tree_5_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var0_source_empty_data;
  reg _add_tree_5_var1_idle;
  reg [33-1:0] _add_tree_5_var1_source_count;
  reg [5-1:0] _add_tree_5_var1_source_mode;
  reg [16-1:0] _add_tree_5_var1_source_generator_id;
  reg [32-1:0] _add_tree_5_var1_source_offset;
  reg [33-1:0] _add_tree_5_var1_source_size;
  reg [32-1:0] _add_tree_5_var1_source_stride;
  reg [32-1:0] _add_tree_5_var1_source_offset_buf;
  reg [33-1:0] _add_tree_5_var1_source_size_buf;
  reg [32-1:0] _add_tree_5_var1_source_stride_buf;
  reg [8-1:0] _add_tree_5_var1_source_sel;
  reg [32-1:0] _add_tree_5_var1_source_ram_raddr;
  reg _add_tree_5_var1_source_ram_renable;
  wire [64-1:0] _add_tree_5_var1_source_ram_rdata;
  reg _add_tree_5_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var1_source_empty_data;
  reg _add_tree_5_var2_idle;
  reg [33-1:0] _add_tree_5_var2_source_count;
  reg [5-1:0] _add_tree_5_var2_source_mode;
  reg [16-1:0] _add_tree_5_var2_source_generator_id;
  reg [32-1:0] _add_tree_5_var2_source_offset;
  reg [33-1:0] _add_tree_5_var2_source_size;
  reg [32-1:0] _add_tree_5_var2_source_stride;
  reg [32-1:0] _add_tree_5_var2_source_offset_buf;
  reg [33-1:0] _add_tree_5_var2_source_size_buf;
  reg [32-1:0] _add_tree_5_var2_source_stride_buf;
  reg [8-1:0] _add_tree_5_var2_source_sel;
  reg [32-1:0] _add_tree_5_var2_source_ram_raddr;
  reg _add_tree_5_var2_source_ram_renable;
  wire [64-1:0] _add_tree_5_var2_source_ram_rdata;
  reg _add_tree_5_var2_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var2_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var2_source_empty_data;
  reg _add_tree_5_var3_idle;
  reg [33-1:0] _add_tree_5_var3_source_count;
  reg [5-1:0] _add_tree_5_var3_source_mode;
  reg [16-1:0] _add_tree_5_var3_source_generator_id;
  reg [32-1:0] _add_tree_5_var3_source_offset;
  reg [33-1:0] _add_tree_5_var3_source_size;
  reg [32-1:0] _add_tree_5_var3_source_stride;
  reg [32-1:0] _add_tree_5_var3_source_offset_buf;
  reg [33-1:0] _add_tree_5_var3_source_size_buf;
  reg [32-1:0] _add_tree_5_var3_source_stride_buf;
  reg [8-1:0] _add_tree_5_var3_source_sel;
  reg [32-1:0] _add_tree_5_var3_source_ram_raddr;
  reg _add_tree_5_var3_source_ram_renable;
  wire [64-1:0] _add_tree_5_var3_source_ram_rdata;
  reg _add_tree_5_var3_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var3_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var3_source_empty_data;
  reg _add_tree_5_var4_idle;
  reg [33-1:0] _add_tree_5_var4_source_count;
  reg [5-1:0] _add_tree_5_var4_source_mode;
  reg [16-1:0] _add_tree_5_var4_source_generator_id;
  reg [32-1:0] _add_tree_5_var4_source_offset;
  reg [33-1:0] _add_tree_5_var4_source_size;
  reg [32-1:0] _add_tree_5_var4_source_stride;
  reg [32-1:0] _add_tree_5_var4_source_offset_buf;
  reg [33-1:0] _add_tree_5_var4_source_size_buf;
  reg [32-1:0] _add_tree_5_var4_source_stride_buf;
  reg [8-1:0] _add_tree_5_var4_source_sel;
  reg [32-1:0] _add_tree_5_var4_source_ram_raddr;
  reg _add_tree_5_var4_source_ram_renable;
  wire [64-1:0] _add_tree_5_var4_source_ram_rdata;
  reg _add_tree_5_var4_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var4_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var4_source_empty_data;
  reg _add_tree_5_var5_idle;
  reg [33-1:0] _add_tree_5_var5_source_count;
  reg [5-1:0] _add_tree_5_var5_source_mode;
  reg [16-1:0] _add_tree_5_var5_source_generator_id;
  reg [32-1:0] _add_tree_5_var5_source_offset;
  reg [33-1:0] _add_tree_5_var5_source_size;
  reg [32-1:0] _add_tree_5_var5_source_stride;
  reg [32-1:0] _add_tree_5_var5_source_offset_buf;
  reg [33-1:0] _add_tree_5_var5_source_size_buf;
  reg [32-1:0] _add_tree_5_var5_source_stride_buf;
  reg [8-1:0] _add_tree_5_var5_source_sel;
  reg [32-1:0] _add_tree_5_var5_source_ram_raddr;
  reg _add_tree_5_var5_source_ram_renable;
  wire [64-1:0] _add_tree_5_var5_source_ram_rdata;
  reg _add_tree_5_var5_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var5_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var5_source_empty_data;
  reg _add_tree_5_var6_idle;
  reg [33-1:0] _add_tree_5_var6_source_count;
  reg [5-1:0] _add_tree_5_var6_source_mode;
  reg [16-1:0] _add_tree_5_var6_source_generator_id;
  reg [32-1:0] _add_tree_5_var6_source_offset;
  reg [33-1:0] _add_tree_5_var6_source_size;
  reg [32-1:0] _add_tree_5_var6_source_stride;
  reg [32-1:0] _add_tree_5_var6_source_offset_buf;
  reg [33-1:0] _add_tree_5_var6_source_size_buf;
  reg [32-1:0] _add_tree_5_var6_source_stride_buf;
  reg [8-1:0] _add_tree_5_var6_source_sel;
  reg [32-1:0] _add_tree_5_var6_source_ram_raddr;
  reg _add_tree_5_var6_source_ram_renable;
  wire [64-1:0] _add_tree_5_var6_source_ram_rdata;
  reg _add_tree_5_var6_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var6_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var6_source_empty_data;
  reg _add_tree_5_var7_idle;
  reg [33-1:0] _add_tree_5_var7_source_count;
  reg [5-1:0] _add_tree_5_var7_source_mode;
  reg [16-1:0] _add_tree_5_var7_source_generator_id;
  reg [32-1:0] _add_tree_5_var7_source_offset;
  reg [33-1:0] _add_tree_5_var7_source_size;
  reg [32-1:0] _add_tree_5_var7_source_stride;
  reg [32-1:0] _add_tree_5_var7_source_offset_buf;
  reg [33-1:0] _add_tree_5_var7_source_size_buf;
  reg [32-1:0] _add_tree_5_var7_source_stride_buf;
  reg [8-1:0] _add_tree_5_var7_source_sel;
  reg [32-1:0] _add_tree_5_var7_source_ram_raddr;
  reg _add_tree_5_var7_source_ram_renable;
  wire [64-1:0] _add_tree_5_var7_source_ram_rdata;
  reg _add_tree_5_var7_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var7_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var7_source_empty_data;
  reg _add_tree_5_var8_idle;
  reg [33-1:0] _add_tree_5_var8_source_count;
  reg [5-1:0] _add_tree_5_var8_source_mode;
  reg [16-1:0] _add_tree_5_var8_source_generator_id;
  reg [32-1:0] _add_tree_5_var8_source_offset;
  reg [33-1:0] _add_tree_5_var8_source_size;
  reg [32-1:0] _add_tree_5_var8_source_stride;
  reg [32-1:0] _add_tree_5_var8_source_offset_buf;
  reg [33-1:0] _add_tree_5_var8_source_size_buf;
  reg [32-1:0] _add_tree_5_var8_source_stride_buf;
  reg [8-1:0] _add_tree_5_var8_source_sel;
  reg [32-1:0] _add_tree_5_var8_source_ram_raddr;
  reg _add_tree_5_var8_source_ram_renable;
  wire [64-1:0] _add_tree_5_var8_source_ram_rdata;
  reg _add_tree_5_var8_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var8_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var8_source_empty_data;
  reg _add_tree_5_var9_idle;
  reg [33-1:0] _add_tree_5_var9_source_count;
  reg [5-1:0] _add_tree_5_var9_source_mode;
  reg [16-1:0] _add_tree_5_var9_source_generator_id;
  reg [32-1:0] _add_tree_5_var9_source_offset;
  reg [33-1:0] _add_tree_5_var9_source_size;
  reg [32-1:0] _add_tree_5_var9_source_stride;
  reg [32-1:0] _add_tree_5_var9_source_offset_buf;
  reg [33-1:0] _add_tree_5_var9_source_size_buf;
  reg [32-1:0] _add_tree_5_var9_source_stride_buf;
  reg [8-1:0] _add_tree_5_var9_source_sel;
  reg [32-1:0] _add_tree_5_var9_source_ram_raddr;
  reg _add_tree_5_var9_source_ram_renable;
  wire [64-1:0] _add_tree_5_var9_source_ram_rdata;
  reg _add_tree_5_var9_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var9_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var9_source_empty_data;
  reg _add_tree_5_var10_idle;
  reg [33-1:0] _add_tree_5_var10_source_count;
  reg [5-1:0] _add_tree_5_var10_source_mode;
  reg [16-1:0] _add_tree_5_var10_source_generator_id;
  reg [32-1:0] _add_tree_5_var10_source_offset;
  reg [33-1:0] _add_tree_5_var10_source_size;
  reg [32-1:0] _add_tree_5_var10_source_stride;
  reg [32-1:0] _add_tree_5_var10_source_offset_buf;
  reg [33-1:0] _add_tree_5_var10_source_size_buf;
  reg [32-1:0] _add_tree_5_var10_source_stride_buf;
  reg [8-1:0] _add_tree_5_var10_source_sel;
  reg [32-1:0] _add_tree_5_var10_source_ram_raddr;
  reg _add_tree_5_var10_source_ram_renable;
  wire [64-1:0] _add_tree_5_var10_source_ram_rdata;
  reg _add_tree_5_var10_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var10_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var10_source_empty_data;
  reg _add_tree_5_var11_idle;
  reg [33-1:0] _add_tree_5_var11_source_count;
  reg [5-1:0] _add_tree_5_var11_source_mode;
  reg [16-1:0] _add_tree_5_var11_source_generator_id;
  reg [32-1:0] _add_tree_5_var11_source_offset;
  reg [33-1:0] _add_tree_5_var11_source_size;
  reg [32-1:0] _add_tree_5_var11_source_stride;
  reg [32-1:0] _add_tree_5_var11_source_offset_buf;
  reg [33-1:0] _add_tree_5_var11_source_size_buf;
  reg [32-1:0] _add_tree_5_var11_source_stride_buf;
  reg [8-1:0] _add_tree_5_var11_source_sel;
  reg [32-1:0] _add_tree_5_var11_source_ram_raddr;
  reg _add_tree_5_var11_source_ram_renable;
  wire [64-1:0] _add_tree_5_var11_source_ram_rdata;
  reg _add_tree_5_var11_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var11_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var11_source_empty_data;
  reg _add_tree_5_var12_idle;
  reg [33-1:0] _add_tree_5_var12_source_count;
  reg [5-1:0] _add_tree_5_var12_source_mode;
  reg [16-1:0] _add_tree_5_var12_source_generator_id;
  reg [32-1:0] _add_tree_5_var12_source_offset;
  reg [33-1:0] _add_tree_5_var12_source_size;
  reg [32-1:0] _add_tree_5_var12_source_stride;
  reg [32-1:0] _add_tree_5_var12_source_offset_buf;
  reg [33-1:0] _add_tree_5_var12_source_size_buf;
  reg [32-1:0] _add_tree_5_var12_source_stride_buf;
  reg [8-1:0] _add_tree_5_var12_source_sel;
  reg [32-1:0] _add_tree_5_var12_source_ram_raddr;
  reg _add_tree_5_var12_source_ram_renable;
  wire [64-1:0] _add_tree_5_var12_source_ram_rdata;
  reg _add_tree_5_var12_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var12_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var12_source_empty_data;
  reg _add_tree_5_var13_idle;
  reg [33-1:0] _add_tree_5_var13_source_count;
  reg [5-1:0] _add_tree_5_var13_source_mode;
  reg [16-1:0] _add_tree_5_var13_source_generator_id;
  reg [32-1:0] _add_tree_5_var13_source_offset;
  reg [33-1:0] _add_tree_5_var13_source_size;
  reg [32-1:0] _add_tree_5_var13_source_stride;
  reg [32-1:0] _add_tree_5_var13_source_offset_buf;
  reg [33-1:0] _add_tree_5_var13_source_size_buf;
  reg [32-1:0] _add_tree_5_var13_source_stride_buf;
  reg [8-1:0] _add_tree_5_var13_source_sel;
  reg [32-1:0] _add_tree_5_var13_source_ram_raddr;
  reg _add_tree_5_var13_source_ram_renable;
  wire [64-1:0] _add_tree_5_var13_source_ram_rdata;
  reg _add_tree_5_var13_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var13_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var13_source_empty_data;
  reg _add_tree_5_var14_idle;
  reg [33-1:0] _add_tree_5_var14_source_count;
  reg [5-1:0] _add_tree_5_var14_source_mode;
  reg [16-1:0] _add_tree_5_var14_source_generator_id;
  reg [32-1:0] _add_tree_5_var14_source_offset;
  reg [33-1:0] _add_tree_5_var14_source_size;
  reg [32-1:0] _add_tree_5_var14_source_stride;
  reg [32-1:0] _add_tree_5_var14_source_offset_buf;
  reg [33-1:0] _add_tree_5_var14_source_size_buf;
  reg [32-1:0] _add_tree_5_var14_source_stride_buf;
  reg [8-1:0] _add_tree_5_var14_source_sel;
  reg [32-1:0] _add_tree_5_var14_source_ram_raddr;
  reg _add_tree_5_var14_source_ram_renable;
  wire [64-1:0] _add_tree_5_var14_source_ram_rdata;
  reg _add_tree_5_var14_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var14_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var14_source_empty_data;
  reg _add_tree_5_var15_idle;
  reg [33-1:0] _add_tree_5_var15_source_count;
  reg [5-1:0] _add_tree_5_var15_source_mode;
  reg [16-1:0] _add_tree_5_var15_source_generator_id;
  reg [32-1:0] _add_tree_5_var15_source_offset;
  reg [33-1:0] _add_tree_5_var15_source_size;
  reg [32-1:0] _add_tree_5_var15_source_stride;
  reg [32-1:0] _add_tree_5_var15_source_offset_buf;
  reg [33-1:0] _add_tree_5_var15_source_size_buf;
  reg [32-1:0] _add_tree_5_var15_source_stride_buf;
  reg [8-1:0] _add_tree_5_var15_source_sel;
  reg [32-1:0] _add_tree_5_var15_source_ram_raddr;
  reg _add_tree_5_var15_source_ram_renable;
  wire [64-1:0] _add_tree_5_var15_source_ram_rdata;
  reg _add_tree_5_var15_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var15_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var15_source_empty_data;
  reg _add_tree_5_var16_idle;
  reg [33-1:0] _add_tree_5_var16_source_count;
  reg [5-1:0] _add_tree_5_var16_source_mode;
  reg [16-1:0] _add_tree_5_var16_source_generator_id;
  reg [32-1:0] _add_tree_5_var16_source_offset;
  reg [33-1:0] _add_tree_5_var16_source_size;
  reg [32-1:0] _add_tree_5_var16_source_stride;
  reg [32-1:0] _add_tree_5_var16_source_offset_buf;
  reg [33-1:0] _add_tree_5_var16_source_size_buf;
  reg [32-1:0] _add_tree_5_var16_source_stride_buf;
  reg [8-1:0] _add_tree_5_var16_source_sel;
  reg [32-1:0] _add_tree_5_var16_source_ram_raddr;
  reg _add_tree_5_var16_source_ram_renable;
  wire [64-1:0] _add_tree_5_var16_source_ram_rdata;
  reg _add_tree_5_var16_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var16_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var16_source_empty_data;
  reg _add_tree_5_var17_idle;
  reg [33-1:0] _add_tree_5_var17_source_count;
  reg [5-1:0] _add_tree_5_var17_source_mode;
  reg [16-1:0] _add_tree_5_var17_source_generator_id;
  reg [32-1:0] _add_tree_5_var17_source_offset;
  reg [33-1:0] _add_tree_5_var17_source_size;
  reg [32-1:0] _add_tree_5_var17_source_stride;
  reg [32-1:0] _add_tree_5_var17_source_offset_buf;
  reg [33-1:0] _add_tree_5_var17_source_size_buf;
  reg [32-1:0] _add_tree_5_var17_source_stride_buf;
  reg [8-1:0] _add_tree_5_var17_source_sel;
  reg [32-1:0] _add_tree_5_var17_source_ram_raddr;
  reg _add_tree_5_var17_source_ram_renable;
  wire [64-1:0] _add_tree_5_var17_source_ram_rdata;
  reg _add_tree_5_var17_source_fifo_deq;
  wire [64-1:0] _add_tree_5_var17_source_fifo_rdata;
  reg [64-1:0] _add_tree_5_var17_source_empty_data;
  reg [33-1:0] _add_tree_5_sum_sink_count;
  reg [5-1:0] _add_tree_5_sum_sink_mode;
  reg [16-1:0] _add_tree_5_sum_sink_generator_id;
  reg [32-1:0] _add_tree_5_sum_sink_offset;
  reg [33-1:0] _add_tree_5_sum_sink_size;
  reg [32-1:0] _add_tree_5_sum_sink_stride;
  reg [32-1:0] _add_tree_5_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_5_sum_sink_size_buf;
  reg [32-1:0] _add_tree_5_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_5_sum_sink_sel;
  reg [32-1:0] _add_tree_5_sum_sink_waddr;
  reg _add_tree_5_sum_sink_wenable;
  reg [64-1:0] _add_tree_5_sum_sink_wdata;
  reg _add_tree_5_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_5_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_5_sum_sink_immediate;
  reg _mul_rshift_round_clip_6_stream_ivalid;
  wire _mul_rshift_round_clip_6_stream_oready;
  wire _mul_rshift_round_clip_6_stream_internal_oready;
  assign _mul_rshift_round_clip_6_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_6_fsm;
  localparam _mul_rshift_round_clip_6_fsm_init = 0;
  wire _mul_rshift_round_clip_6_run_flag;
  assign _mul_rshift_round_clip_6_run_flag = 0;
  reg _mul_rshift_round_clip_6_source_start;
  wire _mul_rshift_round_clip_6_source_stop;
  reg _mul_rshift_round_clip_6_source_busy;
  wire _mul_rshift_round_clip_6_sink_start;
  wire _mul_rshift_round_clip_6_sink_stop;
  wire _mul_rshift_round_clip_6_sink_busy;
  wire _mul_rshift_round_clip_6_busy;
  reg _mul_rshift_round_clip_6_busy_reg;
  wire _mul_rshift_round_clip_6_is_root;
  reg _mul_rshift_round_clip_6_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_6_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_6_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_x_source_ram_raddr;
  reg _mul_rshift_round_clip_6_x_source_ram_renable;
  wire [64-1:0] _mul_rshift_round_clip_6_x_source_ram_rdata;
  reg _mul_rshift_round_clip_6_x_source_fifo_deq;
  wire [64-1:0] _mul_rshift_round_clip_6_x_source_fifo_rdata;
  reg [64-1:0] _mul_rshift_round_clip_6_x_source_empty_data;
  reg _mul_rshift_round_clip_6_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_6_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_6_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_y_source_ram_raddr;
  reg _mul_rshift_round_clip_6_y_source_ram_renable;
  wire [16-1:0] _mul_rshift_round_clip_6_y_source_ram_rdata;
  reg _mul_rshift_round_clip_6_y_source_fifo_deq;
  wire [16-1:0] _mul_rshift_round_clip_6_y_source_fifo_rdata;
  reg [16-1:0] _mul_rshift_round_clip_6_y_source_empty_data;
  reg _mul_rshift_round_clip_6_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_6_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_6_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_6_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_6_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_6_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_6_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_6_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_6_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_6_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_6_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_6_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_6_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_6_z_sink_waddr;
  reg _mul_rshift_round_clip_6_z_sink_wenable;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_wdata;
  reg _mul_rshift_round_clip_6_z_sink_fifo_enq;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_fifo_wdata;
  reg [16-1:0] _mul_rshift_round_clip_6_z_sink_immediate;
  reg _mul_rshift_round_clip_7_stream_ivalid;
  wire _mul_rshift_round_clip_7_stream_oready;
  wire _mul_rshift_round_clip_7_stream_internal_oready;
  assign _mul_rshift_round_clip_7_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_7_fsm;
  localparam _mul_rshift_round_clip_7_fsm_init = 0;
  wire _mul_rshift_round_clip_7_run_flag;
  assign _mul_rshift_round_clip_7_run_flag = 0;
  reg _mul_rshift_round_clip_7_source_start;
  wire _mul_rshift_round_clip_7_source_stop;
  reg _mul_rshift_round_clip_7_source_busy;
  wire _mul_rshift_round_clip_7_sink_start;
  wire _mul_rshift_round_clip_7_sink_stop;
  wire _mul_rshift_round_clip_7_sink_busy;
  wire _mul_rshift_round_clip_7_busy;
  reg _mul_rshift_round_clip_7_busy_reg;
  wire _mul_rshift_round_clip_7_is_root;
  reg _mul_rshift_round_clip_7_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_7_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_7_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_x_source_ram_raddr;
  reg _mul_rshift_round_clip_7_x_source_ram_renable;
  wire [64-1:0] _mul_rshift_round_clip_7_x_source_ram_rdata;
  reg _mul_rshift_round_clip_7_x_source_fifo_deq;
  wire [64-1:0] _mul_rshift_round_clip_7_x_source_fifo_rdata;
  reg [64-1:0] _mul_rshift_round_clip_7_x_source_empty_data;
  reg _mul_rshift_round_clip_7_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_7_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_7_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_y_source_ram_raddr;
  reg _mul_rshift_round_clip_7_y_source_ram_renable;
  wire [16-1:0] _mul_rshift_round_clip_7_y_source_ram_rdata;
  reg _mul_rshift_round_clip_7_y_source_fifo_deq;
  wire [16-1:0] _mul_rshift_round_clip_7_y_source_fifo_rdata;
  reg [16-1:0] _mul_rshift_round_clip_7_y_source_empty_data;
  reg _mul_rshift_round_clip_7_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_7_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_7_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_7_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_7_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_7_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_7_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_7_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_7_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_7_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_7_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_7_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_7_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_7_z_sink_waddr;
  reg _mul_rshift_round_clip_7_z_sink_wenable;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_wdata;
  reg _mul_rshift_round_clip_7_z_sink_fifo_enq;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_fifo_wdata;
  reg [16-1:0] _mul_rshift_round_clip_7_z_sink_immediate;
  reg _mul_8_stream_ivalid;
  wire _mul_8_stream_oready;
  wire _mul_8_stream_internal_oready;
  assign _mul_8_stream_internal_oready = 1;
  reg [32-1:0] _mul_8_fsm;
  localparam _mul_8_fsm_init = 0;
  wire _mul_8_run_flag;
  assign _mul_8_run_flag = 0;
  reg _mul_8_source_start;
  wire _mul_8_source_stop;
  reg _mul_8_source_busy;
  wire _mul_8_sink_start;
  wire _mul_8_sink_stop;
  wire _mul_8_sink_busy;
  wire _mul_8_busy;
  reg _mul_8_busy_reg;
  wire _mul_8_is_root;
  reg _mul_8_x_idle;
  reg [33-1:0] _mul_8_x_source_count;
  reg [5-1:0] _mul_8_x_source_mode;
  reg [16-1:0] _mul_8_x_source_generator_id;
  reg [32-1:0] _mul_8_x_source_offset;
  reg [33-1:0] _mul_8_x_source_size;
  reg [32-1:0] _mul_8_x_source_stride;
  reg [32-1:0] _mul_8_x_source_offset_buf;
  reg [33-1:0] _mul_8_x_source_size_buf;
  reg [32-1:0] _mul_8_x_source_stride_buf;
  reg [8-1:0] _mul_8_x_source_sel;
  reg [32-1:0] _mul_8_x_source_ram_raddr;
  reg _mul_8_x_source_ram_renable;
  wire [16-1:0] _mul_8_x_source_ram_rdata;
  reg _mul_8_x_source_fifo_deq;
  wire [16-1:0] _mul_8_x_source_fifo_rdata;
  reg [16-1:0] _mul_8_x_source_empty_data;
  reg _mul_8_y_idle;
  reg [33-1:0] _mul_8_y_source_count;
  reg [5-1:0] _mul_8_y_source_mode;
  reg [16-1:0] _mul_8_y_source_generator_id;
  reg [32-1:0] _mul_8_y_source_offset;
  reg [33-1:0] _mul_8_y_source_size;
  reg [32-1:0] _mul_8_y_source_stride;
  reg [32-1:0] _mul_8_y_source_offset_buf;
  reg [33-1:0] _mul_8_y_source_size_buf;
  reg [32-1:0] _mul_8_y_source_stride_buf;
  reg [8-1:0] _mul_8_y_source_sel;
  reg [32-1:0] _mul_8_y_source_ram_raddr;
  reg _mul_8_y_source_ram_renable;
  wire [16-1:0] _mul_8_y_source_ram_rdata;
  reg _mul_8_y_source_fifo_deq;
  wire [16-1:0] _mul_8_y_source_fifo_rdata;
  reg [16-1:0] _mul_8_y_source_empty_data;
  reg _mul_8_rshift_idle;
  reg [33-1:0] _mul_8_rshift_source_count;
  reg [5-1:0] _mul_8_rshift_source_mode;
  reg [16-1:0] _mul_8_rshift_source_generator_id;
  reg [32-1:0] _mul_8_rshift_source_offset;
  reg [33-1:0] _mul_8_rshift_source_size;
  reg [32-1:0] _mul_8_rshift_source_stride;
  reg [32-1:0] _mul_8_rshift_source_offset_buf;
  reg [33-1:0] _mul_8_rshift_source_size_buf;
  reg [32-1:0] _mul_8_rshift_source_stride_buf;
  reg [8-1:0] _mul_8_rshift_source_sel;
  reg [32-1:0] _mul_8_rshift_source_ram_raddr;
  reg _mul_8_rshift_source_ram_renable;
  wire [32-1:0] _mul_8_rshift_source_ram_rdata;
  reg _mul_8_rshift_source_fifo_deq;
  wire [32-1:0] _mul_8_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_8_rshift_source_empty_data;
  reg [33-1:0] _mul_8_z_sink_count;
  reg [5-1:0] _mul_8_z_sink_mode;
  reg [16-1:0] _mul_8_z_sink_generator_id;
  reg [32-1:0] _mul_8_z_sink_offset;
  reg [33-1:0] _mul_8_z_sink_size;
  reg [32-1:0] _mul_8_z_sink_stride;
  reg [32-1:0] _mul_8_z_sink_offset_buf;
  reg [33-1:0] _mul_8_z_sink_size_buf;
  reg [32-1:0] _mul_8_z_sink_stride_buf;
  reg [8-1:0] _mul_8_z_sink_sel;
  reg [32-1:0] _mul_8_z_sink_waddr;
  reg _mul_8_z_sink_wenable;
  reg [32-1:0] _mul_8_z_sink_wdata;
  reg _mul_8_z_sink_fifo_enq;
  reg [32-1:0] _mul_8_z_sink_fifo_wdata;
  reg [32-1:0] _mul_8_z_sink_immediate;
  reg _mul_9_stream_ivalid;
  wire _mul_9_stream_oready;
  wire _mul_9_stream_internal_oready;
  assign _mul_9_stream_internal_oready = 1;
  reg [32-1:0] _mul_9_fsm;
  localparam _mul_9_fsm_init = 0;
  wire _mul_9_run_flag;
  assign _mul_9_run_flag = 0;
  reg _mul_9_source_start;
  wire _mul_9_source_stop;
  reg _mul_9_source_busy;
  wire _mul_9_sink_start;
  wire _mul_9_sink_stop;
  wire _mul_9_sink_busy;
  wire _mul_9_busy;
  reg _mul_9_busy_reg;
  wire _mul_9_is_root;
  reg _mul_9_x_idle;
  reg [33-1:0] _mul_9_x_source_count;
  reg [5-1:0] _mul_9_x_source_mode;
  reg [16-1:0] _mul_9_x_source_generator_id;
  reg [32-1:0] _mul_9_x_source_offset;
  reg [33-1:0] _mul_9_x_source_size;
  reg [32-1:0] _mul_9_x_source_stride;
  reg [32-1:0] _mul_9_x_source_offset_buf;
  reg [33-1:0] _mul_9_x_source_size_buf;
  reg [32-1:0] _mul_9_x_source_stride_buf;
  reg [8-1:0] _mul_9_x_source_sel;
  reg [32-1:0] _mul_9_x_source_ram_raddr;
  reg _mul_9_x_source_ram_renable;
  wire [16-1:0] _mul_9_x_source_ram_rdata;
  reg _mul_9_x_source_fifo_deq;
  wire [16-1:0] _mul_9_x_source_fifo_rdata;
  reg [16-1:0] _mul_9_x_source_empty_data;
  reg _mul_9_y_idle;
  reg [33-1:0] _mul_9_y_source_count;
  reg [5-1:0] _mul_9_y_source_mode;
  reg [16-1:0] _mul_9_y_source_generator_id;
  reg [32-1:0] _mul_9_y_source_offset;
  reg [33-1:0] _mul_9_y_source_size;
  reg [32-1:0] _mul_9_y_source_stride;
  reg [32-1:0] _mul_9_y_source_offset_buf;
  reg [33-1:0] _mul_9_y_source_size_buf;
  reg [32-1:0] _mul_9_y_source_stride_buf;
  reg [8-1:0] _mul_9_y_source_sel;
  reg [32-1:0] _mul_9_y_source_ram_raddr;
  reg _mul_9_y_source_ram_renable;
  wire [16-1:0] _mul_9_y_source_ram_rdata;
  reg _mul_9_y_source_fifo_deq;
  wire [16-1:0] _mul_9_y_source_fifo_rdata;
  reg [16-1:0] _mul_9_y_source_empty_data;
  reg _mul_9_rshift_idle;
  reg [33-1:0] _mul_9_rshift_source_count;
  reg [5-1:0] _mul_9_rshift_source_mode;
  reg [16-1:0] _mul_9_rshift_source_generator_id;
  reg [32-1:0] _mul_9_rshift_source_offset;
  reg [33-1:0] _mul_9_rshift_source_size;
  reg [32-1:0] _mul_9_rshift_source_stride;
  reg [32-1:0] _mul_9_rshift_source_offset_buf;
  reg [33-1:0] _mul_9_rshift_source_size_buf;
  reg [32-1:0] _mul_9_rshift_source_stride_buf;
  reg [8-1:0] _mul_9_rshift_source_sel;
  reg [32-1:0] _mul_9_rshift_source_ram_raddr;
  reg _mul_9_rshift_source_ram_renable;
  wire [32-1:0] _mul_9_rshift_source_ram_rdata;
  reg _mul_9_rshift_source_fifo_deq;
  wire [32-1:0] _mul_9_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_9_rshift_source_empty_data;
  reg [33-1:0] _mul_9_z_sink_count;
  reg [5-1:0] _mul_9_z_sink_mode;
  reg [16-1:0] _mul_9_z_sink_generator_id;
  reg [32-1:0] _mul_9_z_sink_offset;
  reg [33-1:0] _mul_9_z_sink_size;
  reg [32-1:0] _mul_9_z_sink_stride;
  reg [32-1:0] _mul_9_z_sink_offset_buf;
  reg [33-1:0] _mul_9_z_sink_size_buf;
  reg [32-1:0] _mul_9_z_sink_stride_buf;
  reg [8-1:0] _mul_9_z_sink_sel;
  reg [32-1:0] _mul_9_z_sink_waddr;
  reg _mul_9_z_sink_wenable;
  reg [32-1:0] _mul_9_z_sink_wdata;
  reg _mul_9_z_sink_fifo_enq;
  reg [32-1:0] _mul_9_z_sink_fifo_wdata;
  reg [32-1:0] _mul_9_z_sink_immediate;
  reg _mul_10_stream_ivalid;
  wire _mul_10_stream_oready;
  wire _mul_10_stream_internal_oready;
  assign _mul_10_stream_internal_oready = 1;
  reg [32-1:0] _mul_10_fsm;
  localparam _mul_10_fsm_init = 0;
  wire _mul_10_run_flag;
  assign _mul_10_run_flag = 0;
  reg _mul_10_source_start;
  wire _mul_10_source_stop;
  reg _mul_10_source_busy;
  wire _mul_10_sink_start;
  wire _mul_10_sink_stop;
  wire _mul_10_sink_busy;
  wire _mul_10_busy;
  reg _mul_10_busy_reg;
  wire _mul_10_is_root;
  reg _mul_10_x_idle;
  reg [33-1:0] _mul_10_x_source_count;
  reg [5-1:0] _mul_10_x_source_mode;
  reg [16-1:0] _mul_10_x_source_generator_id;
  reg [32-1:0] _mul_10_x_source_offset;
  reg [33-1:0] _mul_10_x_source_size;
  reg [32-1:0] _mul_10_x_source_stride;
  reg [32-1:0] _mul_10_x_source_offset_buf;
  reg [33-1:0] _mul_10_x_source_size_buf;
  reg [32-1:0] _mul_10_x_source_stride_buf;
  reg [8-1:0] _mul_10_x_source_sel;
  reg [32-1:0] _mul_10_x_source_ram_raddr;
  reg _mul_10_x_source_ram_renable;
  wire [16-1:0] _mul_10_x_source_ram_rdata;
  reg _mul_10_x_source_fifo_deq;
  wire [16-1:0] _mul_10_x_source_fifo_rdata;
  reg [16-1:0] _mul_10_x_source_empty_data;
  reg _mul_10_y_idle;
  reg [33-1:0] _mul_10_y_source_count;
  reg [5-1:0] _mul_10_y_source_mode;
  reg [16-1:0] _mul_10_y_source_generator_id;
  reg [32-1:0] _mul_10_y_source_offset;
  reg [33-1:0] _mul_10_y_source_size;
  reg [32-1:0] _mul_10_y_source_stride;
  reg [32-1:0] _mul_10_y_source_offset_buf;
  reg [33-1:0] _mul_10_y_source_size_buf;
  reg [32-1:0] _mul_10_y_source_stride_buf;
  reg [8-1:0] _mul_10_y_source_sel;
  reg [32-1:0] _mul_10_y_source_ram_raddr;
  reg _mul_10_y_source_ram_renable;
  wire [16-1:0] _mul_10_y_source_ram_rdata;
  reg _mul_10_y_source_fifo_deq;
  wire [16-1:0] _mul_10_y_source_fifo_rdata;
  reg [16-1:0] _mul_10_y_source_empty_data;
  reg _mul_10_rshift_idle;
  reg [33-1:0] _mul_10_rshift_source_count;
  reg [5-1:0] _mul_10_rshift_source_mode;
  reg [16-1:0] _mul_10_rshift_source_generator_id;
  reg [32-1:0] _mul_10_rshift_source_offset;
  reg [33-1:0] _mul_10_rshift_source_size;
  reg [32-1:0] _mul_10_rshift_source_stride;
  reg [32-1:0] _mul_10_rshift_source_offset_buf;
  reg [33-1:0] _mul_10_rshift_source_size_buf;
  reg [32-1:0] _mul_10_rshift_source_stride_buf;
  reg [8-1:0] _mul_10_rshift_source_sel;
  reg [32-1:0] _mul_10_rshift_source_ram_raddr;
  reg _mul_10_rshift_source_ram_renable;
  wire [32-1:0] _mul_10_rshift_source_ram_rdata;
  reg _mul_10_rshift_source_fifo_deq;
  wire [32-1:0] _mul_10_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_10_rshift_source_empty_data;
  reg [33-1:0] _mul_10_z_sink_count;
  reg [5-1:0] _mul_10_z_sink_mode;
  reg [16-1:0] _mul_10_z_sink_generator_id;
  reg [32-1:0] _mul_10_z_sink_offset;
  reg [33-1:0] _mul_10_z_sink_size;
  reg [32-1:0] _mul_10_z_sink_stride;
  reg [32-1:0] _mul_10_z_sink_offset_buf;
  reg [33-1:0] _mul_10_z_sink_size_buf;
  reg [32-1:0] _mul_10_z_sink_stride_buf;
  reg [8-1:0] _mul_10_z_sink_sel;
  reg [32-1:0] _mul_10_z_sink_waddr;
  reg _mul_10_z_sink_wenable;
  reg [32-1:0] _mul_10_z_sink_wdata;
  reg _mul_10_z_sink_fifo_enq;
  reg [32-1:0] _mul_10_z_sink_fifo_wdata;
  reg [32-1:0] _mul_10_z_sink_immediate;
  reg _mul_11_stream_ivalid;
  wire _mul_11_stream_oready;
  wire _mul_11_stream_internal_oready;
  assign _mul_11_stream_internal_oready = 1;
  reg [32-1:0] _mul_11_fsm;
  localparam _mul_11_fsm_init = 0;
  wire _mul_11_run_flag;
  assign _mul_11_run_flag = 0;
  reg _mul_11_source_start;
  wire _mul_11_source_stop;
  reg _mul_11_source_busy;
  wire _mul_11_sink_start;
  wire _mul_11_sink_stop;
  wire _mul_11_sink_busy;
  wire _mul_11_busy;
  reg _mul_11_busy_reg;
  wire _mul_11_is_root;
  reg _mul_11_x_idle;
  reg [33-1:0] _mul_11_x_source_count;
  reg [5-1:0] _mul_11_x_source_mode;
  reg [16-1:0] _mul_11_x_source_generator_id;
  reg [32-1:0] _mul_11_x_source_offset;
  reg [33-1:0] _mul_11_x_source_size;
  reg [32-1:0] _mul_11_x_source_stride;
  reg [32-1:0] _mul_11_x_source_offset_buf;
  reg [33-1:0] _mul_11_x_source_size_buf;
  reg [32-1:0] _mul_11_x_source_stride_buf;
  reg [8-1:0] _mul_11_x_source_sel;
  reg [32-1:0] _mul_11_x_source_ram_raddr;
  reg _mul_11_x_source_ram_renable;
  wire [16-1:0] _mul_11_x_source_ram_rdata;
  reg _mul_11_x_source_fifo_deq;
  wire [16-1:0] _mul_11_x_source_fifo_rdata;
  reg [16-1:0] _mul_11_x_source_empty_data;
  reg _mul_11_y_idle;
  reg [33-1:0] _mul_11_y_source_count;
  reg [5-1:0] _mul_11_y_source_mode;
  reg [16-1:0] _mul_11_y_source_generator_id;
  reg [32-1:0] _mul_11_y_source_offset;
  reg [33-1:0] _mul_11_y_source_size;
  reg [32-1:0] _mul_11_y_source_stride;
  reg [32-1:0] _mul_11_y_source_offset_buf;
  reg [33-1:0] _mul_11_y_source_size_buf;
  reg [32-1:0] _mul_11_y_source_stride_buf;
  reg [8-1:0] _mul_11_y_source_sel;
  reg [32-1:0] _mul_11_y_source_ram_raddr;
  reg _mul_11_y_source_ram_renable;
  wire [16-1:0] _mul_11_y_source_ram_rdata;
  reg _mul_11_y_source_fifo_deq;
  wire [16-1:0] _mul_11_y_source_fifo_rdata;
  reg [16-1:0] _mul_11_y_source_empty_data;
  reg _mul_11_rshift_idle;
  reg [33-1:0] _mul_11_rshift_source_count;
  reg [5-1:0] _mul_11_rshift_source_mode;
  reg [16-1:0] _mul_11_rshift_source_generator_id;
  reg [32-1:0] _mul_11_rshift_source_offset;
  reg [33-1:0] _mul_11_rshift_source_size;
  reg [32-1:0] _mul_11_rshift_source_stride;
  reg [32-1:0] _mul_11_rshift_source_offset_buf;
  reg [33-1:0] _mul_11_rshift_source_size_buf;
  reg [32-1:0] _mul_11_rshift_source_stride_buf;
  reg [8-1:0] _mul_11_rshift_source_sel;
  reg [32-1:0] _mul_11_rshift_source_ram_raddr;
  reg _mul_11_rshift_source_ram_renable;
  wire [32-1:0] _mul_11_rshift_source_ram_rdata;
  reg _mul_11_rshift_source_fifo_deq;
  wire [32-1:0] _mul_11_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_11_rshift_source_empty_data;
  reg [33-1:0] _mul_11_z_sink_count;
  reg [5-1:0] _mul_11_z_sink_mode;
  reg [16-1:0] _mul_11_z_sink_generator_id;
  reg [32-1:0] _mul_11_z_sink_offset;
  reg [33-1:0] _mul_11_z_sink_size;
  reg [32-1:0] _mul_11_z_sink_stride;
  reg [32-1:0] _mul_11_z_sink_offset_buf;
  reg [33-1:0] _mul_11_z_sink_size_buf;
  reg [32-1:0] _mul_11_z_sink_stride_buf;
  reg [8-1:0] _mul_11_z_sink_sel;
  reg [32-1:0] _mul_11_z_sink_waddr;
  reg _mul_11_z_sink_wenable;
  reg [32-1:0] _mul_11_z_sink_wdata;
  reg _mul_11_z_sink_fifo_enq;
  reg [32-1:0] _mul_11_z_sink_fifo_wdata;
  reg [32-1:0] _mul_11_z_sink_immediate;
  reg _mul_12_stream_ivalid;
  wire _mul_12_stream_oready;
  wire _mul_12_stream_internal_oready;
  assign _mul_12_stream_internal_oready = 1;
  reg [32-1:0] _mul_12_fsm;
  localparam _mul_12_fsm_init = 0;
  wire _mul_12_run_flag;
  assign _mul_12_run_flag = 0;
  reg _mul_12_source_start;
  wire _mul_12_source_stop;
  reg _mul_12_source_busy;
  wire _mul_12_sink_start;
  wire _mul_12_sink_stop;
  wire _mul_12_sink_busy;
  wire _mul_12_busy;
  reg _mul_12_busy_reg;
  wire _mul_12_is_root;
  reg _mul_12_x_idle;
  reg [33-1:0] _mul_12_x_source_count;
  reg [5-1:0] _mul_12_x_source_mode;
  reg [16-1:0] _mul_12_x_source_generator_id;
  reg [32-1:0] _mul_12_x_source_offset;
  reg [33-1:0] _mul_12_x_source_size;
  reg [32-1:0] _mul_12_x_source_stride;
  reg [32-1:0] _mul_12_x_source_offset_buf;
  reg [33-1:0] _mul_12_x_source_size_buf;
  reg [32-1:0] _mul_12_x_source_stride_buf;
  reg [8-1:0] _mul_12_x_source_sel;
  reg [32-1:0] _mul_12_x_source_ram_raddr;
  reg _mul_12_x_source_ram_renable;
  wire [16-1:0] _mul_12_x_source_ram_rdata;
  reg _mul_12_x_source_fifo_deq;
  wire [16-1:0] _mul_12_x_source_fifo_rdata;
  reg [16-1:0] _mul_12_x_source_empty_data;
  reg _mul_12_y_idle;
  reg [33-1:0] _mul_12_y_source_count;
  reg [5-1:0] _mul_12_y_source_mode;
  reg [16-1:0] _mul_12_y_source_generator_id;
  reg [32-1:0] _mul_12_y_source_offset;
  reg [33-1:0] _mul_12_y_source_size;
  reg [32-1:0] _mul_12_y_source_stride;
  reg [32-1:0] _mul_12_y_source_offset_buf;
  reg [33-1:0] _mul_12_y_source_size_buf;
  reg [32-1:0] _mul_12_y_source_stride_buf;
  reg [8-1:0] _mul_12_y_source_sel;
  reg [32-1:0] _mul_12_y_source_ram_raddr;
  reg _mul_12_y_source_ram_renable;
  wire [16-1:0] _mul_12_y_source_ram_rdata;
  reg _mul_12_y_source_fifo_deq;
  wire [16-1:0] _mul_12_y_source_fifo_rdata;
  reg [16-1:0] _mul_12_y_source_empty_data;
  reg _mul_12_rshift_idle;
  reg [33-1:0] _mul_12_rshift_source_count;
  reg [5-1:0] _mul_12_rshift_source_mode;
  reg [16-1:0] _mul_12_rshift_source_generator_id;
  reg [32-1:0] _mul_12_rshift_source_offset;
  reg [33-1:0] _mul_12_rshift_source_size;
  reg [32-1:0] _mul_12_rshift_source_stride;
  reg [32-1:0] _mul_12_rshift_source_offset_buf;
  reg [33-1:0] _mul_12_rshift_source_size_buf;
  reg [32-1:0] _mul_12_rshift_source_stride_buf;
  reg [8-1:0] _mul_12_rshift_source_sel;
  reg [32-1:0] _mul_12_rshift_source_ram_raddr;
  reg _mul_12_rshift_source_ram_renable;
  wire [32-1:0] _mul_12_rshift_source_ram_rdata;
  reg _mul_12_rshift_source_fifo_deq;
  wire [32-1:0] _mul_12_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_12_rshift_source_empty_data;
  reg [33-1:0] _mul_12_z_sink_count;
  reg [5-1:0] _mul_12_z_sink_mode;
  reg [16-1:0] _mul_12_z_sink_generator_id;
  reg [32-1:0] _mul_12_z_sink_offset;
  reg [33-1:0] _mul_12_z_sink_size;
  reg [32-1:0] _mul_12_z_sink_stride;
  reg [32-1:0] _mul_12_z_sink_offset_buf;
  reg [33-1:0] _mul_12_z_sink_size_buf;
  reg [32-1:0] _mul_12_z_sink_stride_buf;
  reg [8-1:0] _mul_12_z_sink_sel;
  reg [32-1:0] _mul_12_z_sink_waddr;
  reg _mul_12_z_sink_wenable;
  reg [32-1:0] _mul_12_z_sink_wdata;
  reg _mul_12_z_sink_fifo_enq;
  reg [32-1:0] _mul_12_z_sink_fifo_wdata;
  reg [32-1:0] _mul_12_z_sink_immediate;
  reg _mul_13_stream_ivalid;
  wire _mul_13_stream_oready;
  wire _mul_13_stream_internal_oready;
  assign _mul_13_stream_internal_oready = 1;
  reg [32-1:0] _mul_13_fsm;
  localparam _mul_13_fsm_init = 0;
  wire _mul_13_run_flag;
  assign _mul_13_run_flag = 0;
  reg _mul_13_source_start;
  wire _mul_13_source_stop;
  reg _mul_13_source_busy;
  wire _mul_13_sink_start;
  wire _mul_13_sink_stop;
  wire _mul_13_sink_busy;
  wire _mul_13_busy;
  reg _mul_13_busy_reg;
  wire _mul_13_is_root;
  reg _mul_13_x_idle;
  reg [33-1:0] _mul_13_x_source_count;
  reg [5-1:0] _mul_13_x_source_mode;
  reg [16-1:0] _mul_13_x_source_generator_id;
  reg [32-1:0] _mul_13_x_source_offset;
  reg [33-1:0] _mul_13_x_source_size;
  reg [32-1:0] _mul_13_x_source_stride;
  reg [32-1:0] _mul_13_x_source_offset_buf;
  reg [33-1:0] _mul_13_x_source_size_buf;
  reg [32-1:0] _mul_13_x_source_stride_buf;
  reg [8-1:0] _mul_13_x_source_sel;
  reg [32-1:0] _mul_13_x_source_ram_raddr;
  reg _mul_13_x_source_ram_renable;
  wire [16-1:0] _mul_13_x_source_ram_rdata;
  reg _mul_13_x_source_fifo_deq;
  wire [16-1:0] _mul_13_x_source_fifo_rdata;
  reg [16-1:0] _mul_13_x_source_empty_data;
  reg _mul_13_y_idle;
  reg [33-1:0] _mul_13_y_source_count;
  reg [5-1:0] _mul_13_y_source_mode;
  reg [16-1:0] _mul_13_y_source_generator_id;
  reg [32-1:0] _mul_13_y_source_offset;
  reg [33-1:0] _mul_13_y_source_size;
  reg [32-1:0] _mul_13_y_source_stride;
  reg [32-1:0] _mul_13_y_source_offset_buf;
  reg [33-1:0] _mul_13_y_source_size_buf;
  reg [32-1:0] _mul_13_y_source_stride_buf;
  reg [8-1:0] _mul_13_y_source_sel;
  reg [32-1:0] _mul_13_y_source_ram_raddr;
  reg _mul_13_y_source_ram_renable;
  wire [16-1:0] _mul_13_y_source_ram_rdata;
  reg _mul_13_y_source_fifo_deq;
  wire [16-1:0] _mul_13_y_source_fifo_rdata;
  reg [16-1:0] _mul_13_y_source_empty_data;
  reg _mul_13_rshift_idle;
  reg [33-1:0] _mul_13_rshift_source_count;
  reg [5-1:0] _mul_13_rshift_source_mode;
  reg [16-1:0] _mul_13_rshift_source_generator_id;
  reg [32-1:0] _mul_13_rshift_source_offset;
  reg [33-1:0] _mul_13_rshift_source_size;
  reg [32-1:0] _mul_13_rshift_source_stride;
  reg [32-1:0] _mul_13_rshift_source_offset_buf;
  reg [33-1:0] _mul_13_rshift_source_size_buf;
  reg [32-1:0] _mul_13_rshift_source_stride_buf;
  reg [8-1:0] _mul_13_rshift_source_sel;
  reg [32-1:0] _mul_13_rshift_source_ram_raddr;
  reg _mul_13_rshift_source_ram_renable;
  wire [32-1:0] _mul_13_rshift_source_ram_rdata;
  reg _mul_13_rshift_source_fifo_deq;
  wire [32-1:0] _mul_13_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_13_rshift_source_empty_data;
  reg [33-1:0] _mul_13_z_sink_count;
  reg [5-1:0] _mul_13_z_sink_mode;
  reg [16-1:0] _mul_13_z_sink_generator_id;
  reg [32-1:0] _mul_13_z_sink_offset;
  reg [33-1:0] _mul_13_z_sink_size;
  reg [32-1:0] _mul_13_z_sink_stride;
  reg [32-1:0] _mul_13_z_sink_offset_buf;
  reg [33-1:0] _mul_13_z_sink_size_buf;
  reg [32-1:0] _mul_13_z_sink_stride_buf;
  reg [8-1:0] _mul_13_z_sink_sel;
  reg [32-1:0] _mul_13_z_sink_waddr;
  reg _mul_13_z_sink_wenable;
  reg [32-1:0] _mul_13_z_sink_wdata;
  reg _mul_13_z_sink_fifo_enq;
  reg [32-1:0] _mul_13_z_sink_fifo_wdata;
  reg [32-1:0] _mul_13_z_sink_immediate;
  reg _mul_14_stream_ivalid;
  wire _mul_14_stream_oready;
  wire _mul_14_stream_internal_oready;
  assign _mul_14_stream_internal_oready = 1;
  reg [32-1:0] _mul_14_fsm;
  localparam _mul_14_fsm_init = 0;
  wire _mul_14_run_flag;
  assign _mul_14_run_flag = 0;
  reg _mul_14_source_start;
  wire _mul_14_source_stop;
  reg _mul_14_source_busy;
  wire _mul_14_sink_start;
  wire _mul_14_sink_stop;
  wire _mul_14_sink_busy;
  wire _mul_14_busy;
  reg _mul_14_busy_reg;
  wire _mul_14_is_root;
  reg _mul_14_x_idle;
  reg [33-1:0] _mul_14_x_source_count;
  reg [5-1:0] _mul_14_x_source_mode;
  reg [16-1:0] _mul_14_x_source_generator_id;
  reg [32-1:0] _mul_14_x_source_offset;
  reg [33-1:0] _mul_14_x_source_size;
  reg [32-1:0] _mul_14_x_source_stride;
  reg [32-1:0] _mul_14_x_source_offset_buf;
  reg [33-1:0] _mul_14_x_source_size_buf;
  reg [32-1:0] _mul_14_x_source_stride_buf;
  reg [8-1:0] _mul_14_x_source_sel;
  reg [32-1:0] _mul_14_x_source_ram_raddr;
  reg _mul_14_x_source_ram_renable;
  wire [16-1:0] _mul_14_x_source_ram_rdata;
  reg _mul_14_x_source_fifo_deq;
  wire [16-1:0] _mul_14_x_source_fifo_rdata;
  reg [16-1:0] _mul_14_x_source_empty_data;
  reg _mul_14_y_idle;
  reg [33-1:0] _mul_14_y_source_count;
  reg [5-1:0] _mul_14_y_source_mode;
  reg [16-1:0] _mul_14_y_source_generator_id;
  reg [32-1:0] _mul_14_y_source_offset;
  reg [33-1:0] _mul_14_y_source_size;
  reg [32-1:0] _mul_14_y_source_stride;
  reg [32-1:0] _mul_14_y_source_offset_buf;
  reg [33-1:0] _mul_14_y_source_size_buf;
  reg [32-1:0] _mul_14_y_source_stride_buf;
  reg [8-1:0] _mul_14_y_source_sel;
  reg [32-1:0] _mul_14_y_source_ram_raddr;
  reg _mul_14_y_source_ram_renable;
  wire [16-1:0] _mul_14_y_source_ram_rdata;
  reg _mul_14_y_source_fifo_deq;
  wire [16-1:0] _mul_14_y_source_fifo_rdata;
  reg [16-1:0] _mul_14_y_source_empty_data;
  reg _mul_14_rshift_idle;
  reg [33-1:0] _mul_14_rshift_source_count;
  reg [5-1:0] _mul_14_rshift_source_mode;
  reg [16-1:0] _mul_14_rshift_source_generator_id;
  reg [32-1:0] _mul_14_rshift_source_offset;
  reg [33-1:0] _mul_14_rshift_source_size;
  reg [32-1:0] _mul_14_rshift_source_stride;
  reg [32-1:0] _mul_14_rshift_source_offset_buf;
  reg [33-1:0] _mul_14_rshift_source_size_buf;
  reg [32-1:0] _mul_14_rshift_source_stride_buf;
  reg [8-1:0] _mul_14_rshift_source_sel;
  reg [32-1:0] _mul_14_rshift_source_ram_raddr;
  reg _mul_14_rshift_source_ram_renable;
  wire [32-1:0] _mul_14_rshift_source_ram_rdata;
  reg _mul_14_rshift_source_fifo_deq;
  wire [32-1:0] _mul_14_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_14_rshift_source_empty_data;
  reg [33-1:0] _mul_14_z_sink_count;
  reg [5-1:0] _mul_14_z_sink_mode;
  reg [16-1:0] _mul_14_z_sink_generator_id;
  reg [32-1:0] _mul_14_z_sink_offset;
  reg [33-1:0] _mul_14_z_sink_size;
  reg [32-1:0] _mul_14_z_sink_stride;
  reg [32-1:0] _mul_14_z_sink_offset_buf;
  reg [33-1:0] _mul_14_z_sink_size_buf;
  reg [32-1:0] _mul_14_z_sink_stride_buf;
  reg [8-1:0] _mul_14_z_sink_sel;
  reg [32-1:0] _mul_14_z_sink_waddr;
  reg _mul_14_z_sink_wenable;
  reg [32-1:0] _mul_14_z_sink_wdata;
  reg _mul_14_z_sink_fifo_enq;
  reg [32-1:0] _mul_14_z_sink_fifo_wdata;
  reg [32-1:0] _mul_14_z_sink_immediate;
  reg _mul_15_stream_ivalid;
  wire _mul_15_stream_oready;
  wire _mul_15_stream_internal_oready;
  assign _mul_15_stream_internal_oready = 1;
  reg [32-1:0] _mul_15_fsm;
  localparam _mul_15_fsm_init = 0;
  wire _mul_15_run_flag;
  assign _mul_15_run_flag = 0;
  reg _mul_15_source_start;
  wire _mul_15_source_stop;
  reg _mul_15_source_busy;
  wire _mul_15_sink_start;
  wire _mul_15_sink_stop;
  wire _mul_15_sink_busy;
  wire _mul_15_busy;
  reg _mul_15_busy_reg;
  wire _mul_15_is_root;
  reg _mul_15_x_idle;
  reg [33-1:0] _mul_15_x_source_count;
  reg [5-1:0] _mul_15_x_source_mode;
  reg [16-1:0] _mul_15_x_source_generator_id;
  reg [32-1:0] _mul_15_x_source_offset;
  reg [33-1:0] _mul_15_x_source_size;
  reg [32-1:0] _mul_15_x_source_stride;
  reg [32-1:0] _mul_15_x_source_offset_buf;
  reg [33-1:0] _mul_15_x_source_size_buf;
  reg [32-1:0] _mul_15_x_source_stride_buf;
  reg [8-1:0] _mul_15_x_source_sel;
  reg [32-1:0] _mul_15_x_source_ram_raddr;
  reg _mul_15_x_source_ram_renable;
  wire [16-1:0] _mul_15_x_source_ram_rdata;
  reg _mul_15_x_source_fifo_deq;
  wire [16-1:0] _mul_15_x_source_fifo_rdata;
  reg [16-1:0] _mul_15_x_source_empty_data;
  reg _mul_15_y_idle;
  reg [33-1:0] _mul_15_y_source_count;
  reg [5-1:0] _mul_15_y_source_mode;
  reg [16-1:0] _mul_15_y_source_generator_id;
  reg [32-1:0] _mul_15_y_source_offset;
  reg [33-1:0] _mul_15_y_source_size;
  reg [32-1:0] _mul_15_y_source_stride;
  reg [32-1:0] _mul_15_y_source_offset_buf;
  reg [33-1:0] _mul_15_y_source_size_buf;
  reg [32-1:0] _mul_15_y_source_stride_buf;
  reg [8-1:0] _mul_15_y_source_sel;
  reg [32-1:0] _mul_15_y_source_ram_raddr;
  reg _mul_15_y_source_ram_renable;
  wire [16-1:0] _mul_15_y_source_ram_rdata;
  reg _mul_15_y_source_fifo_deq;
  wire [16-1:0] _mul_15_y_source_fifo_rdata;
  reg [16-1:0] _mul_15_y_source_empty_data;
  reg _mul_15_rshift_idle;
  reg [33-1:0] _mul_15_rshift_source_count;
  reg [5-1:0] _mul_15_rshift_source_mode;
  reg [16-1:0] _mul_15_rshift_source_generator_id;
  reg [32-1:0] _mul_15_rshift_source_offset;
  reg [33-1:0] _mul_15_rshift_source_size;
  reg [32-1:0] _mul_15_rshift_source_stride;
  reg [32-1:0] _mul_15_rshift_source_offset_buf;
  reg [33-1:0] _mul_15_rshift_source_size_buf;
  reg [32-1:0] _mul_15_rshift_source_stride_buf;
  reg [8-1:0] _mul_15_rshift_source_sel;
  reg [32-1:0] _mul_15_rshift_source_ram_raddr;
  reg _mul_15_rshift_source_ram_renable;
  wire [32-1:0] _mul_15_rshift_source_ram_rdata;
  reg _mul_15_rshift_source_fifo_deq;
  wire [32-1:0] _mul_15_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_15_rshift_source_empty_data;
  reg [33-1:0] _mul_15_z_sink_count;
  reg [5-1:0] _mul_15_z_sink_mode;
  reg [16-1:0] _mul_15_z_sink_generator_id;
  reg [32-1:0] _mul_15_z_sink_offset;
  reg [33-1:0] _mul_15_z_sink_size;
  reg [32-1:0] _mul_15_z_sink_stride;
  reg [32-1:0] _mul_15_z_sink_offset_buf;
  reg [33-1:0] _mul_15_z_sink_size_buf;
  reg [32-1:0] _mul_15_z_sink_stride_buf;
  reg [8-1:0] _mul_15_z_sink_sel;
  reg [32-1:0] _mul_15_z_sink_waddr;
  reg _mul_15_z_sink_wenable;
  reg [32-1:0] _mul_15_z_sink_wdata;
  reg _mul_15_z_sink_fifo_enq;
  reg [32-1:0] _mul_15_z_sink_fifo_wdata;
  reg [32-1:0] _mul_15_z_sink_immediate;
  reg _mul_16_stream_ivalid;
  wire _mul_16_stream_oready;
  wire _mul_16_stream_internal_oready;
  assign _mul_16_stream_internal_oready = 1;
  reg [32-1:0] _mul_16_fsm;
  localparam _mul_16_fsm_init = 0;
  wire _mul_16_run_flag;
  assign _mul_16_run_flag = 0;
  reg _mul_16_source_start;
  wire _mul_16_source_stop;
  reg _mul_16_source_busy;
  wire _mul_16_sink_start;
  wire _mul_16_sink_stop;
  wire _mul_16_sink_busy;
  wire _mul_16_busy;
  reg _mul_16_busy_reg;
  wire _mul_16_is_root;
  reg _mul_16_x_idle;
  reg [33-1:0] _mul_16_x_source_count;
  reg [5-1:0] _mul_16_x_source_mode;
  reg [16-1:0] _mul_16_x_source_generator_id;
  reg [32-1:0] _mul_16_x_source_offset;
  reg [33-1:0] _mul_16_x_source_size;
  reg [32-1:0] _mul_16_x_source_stride;
  reg [32-1:0] _mul_16_x_source_offset_buf;
  reg [33-1:0] _mul_16_x_source_size_buf;
  reg [32-1:0] _mul_16_x_source_stride_buf;
  reg [8-1:0] _mul_16_x_source_sel;
  reg [32-1:0] _mul_16_x_source_ram_raddr;
  reg _mul_16_x_source_ram_renable;
  wire [16-1:0] _mul_16_x_source_ram_rdata;
  reg _mul_16_x_source_fifo_deq;
  wire [16-1:0] _mul_16_x_source_fifo_rdata;
  reg [16-1:0] _mul_16_x_source_empty_data;
  reg _mul_16_y_idle;
  reg [33-1:0] _mul_16_y_source_count;
  reg [5-1:0] _mul_16_y_source_mode;
  reg [16-1:0] _mul_16_y_source_generator_id;
  reg [32-1:0] _mul_16_y_source_offset;
  reg [33-1:0] _mul_16_y_source_size;
  reg [32-1:0] _mul_16_y_source_stride;
  reg [32-1:0] _mul_16_y_source_offset_buf;
  reg [33-1:0] _mul_16_y_source_size_buf;
  reg [32-1:0] _mul_16_y_source_stride_buf;
  reg [8-1:0] _mul_16_y_source_sel;
  reg [32-1:0] _mul_16_y_source_ram_raddr;
  reg _mul_16_y_source_ram_renable;
  wire [16-1:0] _mul_16_y_source_ram_rdata;
  reg _mul_16_y_source_fifo_deq;
  wire [16-1:0] _mul_16_y_source_fifo_rdata;
  reg [16-1:0] _mul_16_y_source_empty_data;
  reg _mul_16_rshift_idle;
  reg [33-1:0] _mul_16_rshift_source_count;
  reg [5-1:0] _mul_16_rshift_source_mode;
  reg [16-1:0] _mul_16_rshift_source_generator_id;
  reg [32-1:0] _mul_16_rshift_source_offset;
  reg [33-1:0] _mul_16_rshift_source_size;
  reg [32-1:0] _mul_16_rshift_source_stride;
  reg [32-1:0] _mul_16_rshift_source_offset_buf;
  reg [33-1:0] _mul_16_rshift_source_size_buf;
  reg [32-1:0] _mul_16_rshift_source_stride_buf;
  reg [8-1:0] _mul_16_rshift_source_sel;
  reg [32-1:0] _mul_16_rshift_source_ram_raddr;
  reg _mul_16_rshift_source_ram_renable;
  wire [32-1:0] _mul_16_rshift_source_ram_rdata;
  reg _mul_16_rshift_source_fifo_deq;
  wire [32-1:0] _mul_16_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_16_rshift_source_empty_data;
  reg [33-1:0] _mul_16_z_sink_count;
  reg [5-1:0] _mul_16_z_sink_mode;
  reg [16-1:0] _mul_16_z_sink_generator_id;
  reg [32-1:0] _mul_16_z_sink_offset;
  reg [33-1:0] _mul_16_z_sink_size;
  reg [32-1:0] _mul_16_z_sink_stride;
  reg [32-1:0] _mul_16_z_sink_offset_buf;
  reg [33-1:0] _mul_16_z_sink_size_buf;
  reg [32-1:0] _mul_16_z_sink_stride_buf;
  reg [8-1:0] _mul_16_z_sink_sel;
  reg [32-1:0] _mul_16_z_sink_waddr;
  reg _mul_16_z_sink_wenable;
  reg [32-1:0] _mul_16_z_sink_wdata;
  reg _mul_16_z_sink_fifo_enq;
  reg [32-1:0] _mul_16_z_sink_fifo_wdata;
  reg [32-1:0] _mul_16_z_sink_immediate;
  reg _mul_17_stream_ivalid;
  wire _mul_17_stream_oready;
  wire _mul_17_stream_internal_oready;
  assign _mul_17_stream_internal_oready = 1;
  reg [32-1:0] _mul_17_fsm;
  localparam _mul_17_fsm_init = 0;
  wire _mul_17_run_flag;
  assign _mul_17_run_flag = 0;
  reg _mul_17_source_start;
  wire _mul_17_source_stop;
  reg _mul_17_source_busy;
  wire _mul_17_sink_start;
  wire _mul_17_sink_stop;
  wire _mul_17_sink_busy;
  wire _mul_17_busy;
  reg _mul_17_busy_reg;
  wire _mul_17_is_root;
  reg _mul_17_x_idle;
  reg [33-1:0] _mul_17_x_source_count;
  reg [5-1:0] _mul_17_x_source_mode;
  reg [16-1:0] _mul_17_x_source_generator_id;
  reg [32-1:0] _mul_17_x_source_offset;
  reg [33-1:0] _mul_17_x_source_size;
  reg [32-1:0] _mul_17_x_source_stride;
  reg [32-1:0] _mul_17_x_source_offset_buf;
  reg [33-1:0] _mul_17_x_source_size_buf;
  reg [32-1:0] _mul_17_x_source_stride_buf;
  reg [8-1:0] _mul_17_x_source_sel;
  reg [32-1:0] _mul_17_x_source_ram_raddr;
  reg _mul_17_x_source_ram_renable;
  wire [16-1:0] _mul_17_x_source_ram_rdata;
  reg _mul_17_x_source_fifo_deq;
  wire [16-1:0] _mul_17_x_source_fifo_rdata;
  reg [16-1:0] _mul_17_x_source_empty_data;
  reg _mul_17_y_idle;
  reg [33-1:0] _mul_17_y_source_count;
  reg [5-1:0] _mul_17_y_source_mode;
  reg [16-1:0] _mul_17_y_source_generator_id;
  reg [32-1:0] _mul_17_y_source_offset;
  reg [33-1:0] _mul_17_y_source_size;
  reg [32-1:0] _mul_17_y_source_stride;
  reg [32-1:0] _mul_17_y_source_offset_buf;
  reg [33-1:0] _mul_17_y_source_size_buf;
  reg [32-1:0] _mul_17_y_source_stride_buf;
  reg [8-1:0] _mul_17_y_source_sel;
  reg [32-1:0] _mul_17_y_source_ram_raddr;
  reg _mul_17_y_source_ram_renable;
  wire [16-1:0] _mul_17_y_source_ram_rdata;
  reg _mul_17_y_source_fifo_deq;
  wire [16-1:0] _mul_17_y_source_fifo_rdata;
  reg [16-1:0] _mul_17_y_source_empty_data;
  reg _mul_17_rshift_idle;
  reg [33-1:0] _mul_17_rshift_source_count;
  reg [5-1:0] _mul_17_rshift_source_mode;
  reg [16-1:0] _mul_17_rshift_source_generator_id;
  reg [32-1:0] _mul_17_rshift_source_offset;
  reg [33-1:0] _mul_17_rshift_source_size;
  reg [32-1:0] _mul_17_rshift_source_stride;
  reg [32-1:0] _mul_17_rshift_source_offset_buf;
  reg [33-1:0] _mul_17_rshift_source_size_buf;
  reg [32-1:0] _mul_17_rshift_source_stride_buf;
  reg [8-1:0] _mul_17_rshift_source_sel;
  reg [32-1:0] _mul_17_rshift_source_ram_raddr;
  reg _mul_17_rshift_source_ram_renable;
  wire [32-1:0] _mul_17_rshift_source_ram_rdata;
  reg _mul_17_rshift_source_fifo_deq;
  wire [32-1:0] _mul_17_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_17_rshift_source_empty_data;
  reg [33-1:0] _mul_17_z_sink_count;
  reg [5-1:0] _mul_17_z_sink_mode;
  reg [16-1:0] _mul_17_z_sink_generator_id;
  reg [32-1:0] _mul_17_z_sink_offset;
  reg [33-1:0] _mul_17_z_sink_size;
  reg [32-1:0] _mul_17_z_sink_stride;
  reg [32-1:0] _mul_17_z_sink_offset_buf;
  reg [33-1:0] _mul_17_z_sink_size_buf;
  reg [32-1:0] _mul_17_z_sink_stride_buf;
  reg [8-1:0] _mul_17_z_sink_sel;
  reg [32-1:0] _mul_17_z_sink_waddr;
  reg _mul_17_z_sink_wenable;
  reg [32-1:0] _mul_17_z_sink_wdata;
  reg _mul_17_z_sink_fifo_enq;
  reg [32-1:0] _mul_17_z_sink_fifo_wdata;
  reg [32-1:0] _mul_17_z_sink_immediate;
  reg _mul_18_stream_ivalid;
  wire _mul_18_stream_oready;
  wire _mul_18_stream_internal_oready;
  assign _mul_18_stream_internal_oready = 1;
  reg [32-1:0] _mul_18_fsm;
  localparam _mul_18_fsm_init = 0;
  wire _mul_18_run_flag;
  assign _mul_18_run_flag = 0;
  reg _mul_18_source_start;
  wire _mul_18_source_stop;
  reg _mul_18_source_busy;
  wire _mul_18_sink_start;
  wire _mul_18_sink_stop;
  wire _mul_18_sink_busy;
  wire _mul_18_busy;
  reg _mul_18_busy_reg;
  wire _mul_18_is_root;
  reg _mul_18_x_idle;
  reg [33-1:0] _mul_18_x_source_count;
  reg [5-1:0] _mul_18_x_source_mode;
  reg [16-1:0] _mul_18_x_source_generator_id;
  reg [32-1:0] _mul_18_x_source_offset;
  reg [33-1:0] _mul_18_x_source_size;
  reg [32-1:0] _mul_18_x_source_stride;
  reg [32-1:0] _mul_18_x_source_offset_buf;
  reg [33-1:0] _mul_18_x_source_size_buf;
  reg [32-1:0] _mul_18_x_source_stride_buf;
  reg [8-1:0] _mul_18_x_source_sel;
  reg [32-1:0] _mul_18_x_source_ram_raddr;
  reg _mul_18_x_source_ram_renable;
  wire [16-1:0] _mul_18_x_source_ram_rdata;
  reg _mul_18_x_source_fifo_deq;
  wire [16-1:0] _mul_18_x_source_fifo_rdata;
  reg [16-1:0] _mul_18_x_source_empty_data;
  reg _mul_18_y_idle;
  reg [33-1:0] _mul_18_y_source_count;
  reg [5-1:0] _mul_18_y_source_mode;
  reg [16-1:0] _mul_18_y_source_generator_id;
  reg [32-1:0] _mul_18_y_source_offset;
  reg [33-1:0] _mul_18_y_source_size;
  reg [32-1:0] _mul_18_y_source_stride;
  reg [32-1:0] _mul_18_y_source_offset_buf;
  reg [33-1:0] _mul_18_y_source_size_buf;
  reg [32-1:0] _mul_18_y_source_stride_buf;
  reg [8-1:0] _mul_18_y_source_sel;
  reg [32-1:0] _mul_18_y_source_ram_raddr;
  reg _mul_18_y_source_ram_renable;
  wire [16-1:0] _mul_18_y_source_ram_rdata;
  reg _mul_18_y_source_fifo_deq;
  wire [16-1:0] _mul_18_y_source_fifo_rdata;
  reg [16-1:0] _mul_18_y_source_empty_data;
  reg _mul_18_rshift_idle;
  reg [33-1:0] _mul_18_rshift_source_count;
  reg [5-1:0] _mul_18_rshift_source_mode;
  reg [16-1:0] _mul_18_rshift_source_generator_id;
  reg [32-1:0] _mul_18_rshift_source_offset;
  reg [33-1:0] _mul_18_rshift_source_size;
  reg [32-1:0] _mul_18_rshift_source_stride;
  reg [32-1:0] _mul_18_rshift_source_offset_buf;
  reg [33-1:0] _mul_18_rshift_source_size_buf;
  reg [32-1:0] _mul_18_rshift_source_stride_buf;
  reg [8-1:0] _mul_18_rshift_source_sel;
  reg [32-1:0] _mul_18_rshift_source_ram_raddr;
  reg _mul_18_rshift_source_ram_renable;
  wire [32-1:0] _mul_18_rshift_source_ram_rdata;
  reg _mul_18_rshift_source_fifo_deq;
  wire [32-1:0] _mul_18_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_18_rshift_source_empty_data;
  reg [33-1:0] _mul_18_z_sink_count;
  reg [5-1:0] _mul_18_z_sink_mode;
  reg [16-1:0] _mul_18_z_sink_generator_id;
  reg [32-1:0] _mul_18_z_sink_offset;
  reg [33-1:0] _mul_18_z_sink_size;
  reg [32-1:0] _mul_18_z_sink_stride;
  reg [32-1:0] _mul_18_z_sink_offset_buf;
  reg [33-1:0] _mul_18_z_sink_size_buf;
  reg [32-1:0] _mul_18_z_sink_stride_buf;
  reg [8-1:0] _mul_18_z_sink_sel;
  reg [32-1:0] _mul_18_z_sink_waddr;
  reg _mul_18_z_sink_wenable;
  reg [32-1:0] _mul_18_z_sink_wdata;
  reg _mul_18_z_sink_fifo_enq;
  reg [32-1:0] _mul_18_z_sink_fifo_wdata;
  reg [32-1:0] _mul_18_z_sink_immediate;
  reg _mul_19_stream_ivalid;
  wire _mul_19_stream_oready;
  wire _mul_19_stream_internal_oready;
  assign _mul_19_stream_internal_oready = 1;
  reg [32-1:0] _mul_19_fsm;
  localparam _mul_19_fsm_init = 0;
  wire _mul_19_run_flag;
  assign _mul_19_run_flag = 0;
  reg _mul_19_source_start;
  wire _mul_19_source_stop;
  reg _mul_19_source_busy;
  wire _mul_19_sink_start;
  wire _mul_19_sink_stop;
  wire _mul_19_sink_busy;
  wire _mul_19_busy;
  reg _mul_19_busy_reg;
  wire _mul_19_is_root;
  reg _mul_19_x_idle;
  reg [33-1:0] _mul_19_x_source_count;
  reg [5-1:0] _mul_19_x_source_mode;
  reg [16-1:0] _mul_19_x_source_generator_id;
  reg [32-1:0] _mul_19_x_source_offset;
  reg [33-1:0] _mul_19_x_source_size;
  reg [32-1:0] _mul_19_x_source_stride;
  reg [32-1:0] _mul_19_x_source_offset_buf;
  reg [33-1:0] _mul_19_x_source_size_buf;
  reg [32-1:0] _mul_19_x_source_stride_buf;
  reg [8-1:0] _mul_19_x_source_sel;
  reg [32-1:0] _mul_19_x_source_ram_raddr;
  reg _mul_19_x_source_ram_renable;
  wire [16-1:0] _mul_19_x_source_ram_rdata;
  reg _mul_19_x_source_fifo_deq;
  wire [16-1:0] _mul_19_x_source_fifo_rdata;
  reg [16-1:0] _mul_19_x_source_empty_data;
  reg _mul_19_y_idle;
  reg [33-1:0] _mul_19_y_source_count;
  reg [5-1:0] _mul_19_y_source_mode;
  reg [16-1:0] _mul_19_y_source_generator_id;
  reg [32-1:0] _mul_19_y_source_offset;
  reg [33-1:0] _mul_19_y_source_size;
  reg [32-1:0] _mul_19_y_source_stride;
  reg [32-1:0] _mul_19_y_source_offset_buf;
  reg [33-1:0] _mul_19_y_source_size_buf;
  reg [32-1:0] _mul_19_y_source_stride_buf;
  reg [8-1:0] _mul_19_y_source_sel;
  reg [32-1:0] _mul_19_y_source_ram_raddr;
  reg _mul_19_y_source_ram_renable;
  wire [16-1:0] _mul_19_y_source_ram_rdata;
  reg _mul_19_y_source_fifo_deq;
  wire [16-1:0] _mul_19_y_source_fifo_rdata;
  reg [16-1:0] _mul_19_y_source_empty_data;
  reg _mul_19_rshift_idle;
  reg [33-1:0] _mul_19_rshift_source_count;
  reg [5-1:0] _mul_19_rshift_source_mode;
  reg [16-1:0] _mul_19_rshift_source_generator_id;
  reg [32-1:0] _mul_19_rshift_source_offset;
  reg [33-1:0] _mul_19_rshift_source_size;
  reg [32-1:0] _mul_19_rshift_source_stride;
  reg [32-1:0] _mul_19_rshift_source_offset_buf;
  reg [33-1:0] _mul_19_rshift_source_size_buf;
  reg [32-1:0] _mul_19_rshift_source_stride_buf;
  reg [8-1:0] _mul_19_rshift_source_sel;
  reg [32-1:0] _mul_19_rshift_source_ram_raddr;
  reg _mul_19_rshift_source_ram_renable;
  wire [32-1:0] _mul_19_rshift_source_ram_rdata;
  reg _mul_19_rshift_source_fifo_deq;
  wire [32-1:0] _mul_19_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_19_rshift_source_empty_data;
  reg [33-1:0] _mul_19_z_sink_count;
  reg [5-1:0] _mul_19_z_sink_mode;
  reg [16-1:0] _mul_19_z_sink_generator_id;
  reg [32-1:0] _mul_19_z_sink_offset;
  reg [33-1:0] _mul_19_z_sink_size;
  reg [32-1:0] _mul_19_z_sink_stride;
  reg [32-1:0] _mul_19_z_sink_offset_buf;
  reg [33-1:0] _mul_19_z_sink_size_buf;
  reg [32-1:0] _mul_19_z_sink_stride_buf;
  reg [8-1:0] _mul_19_z_sink_sel;
  reg [32-1:0] _mul_19_z_sink_waddr;
  reg _mul_19_z_sink_wenable;
  reg [32-1:0] _mul_19_z_sink_wdata;
  reg _mul_19_z_sink_fifo_enq;
  reg [32-1:0] _mul_19_z_sink_fifo_wdata;
  reg [32-1:0] _mul_19_z_sink_immediate;
  reg _mul_20_stream_ivalid;
  wire _mul_20_stream_oready;
  wire _mul_20_stream_internal_oready;
  assign _mul_20_stream_internal_oready = 1;
  reg [32-1:0] _mul_20_fsm;
  localparam _mul_20_fsm_init = 0;
  wire _mul_20_run_flag;
  assign _mul_20_run_flag = 0;
  reg _mul_20_source_start;
  wire _mul_20_source_stop;
  reg _mul_20_source_busy;
  wire _mul_20_sink_start;
  wire _mul_20_sink_stop;
  wire _mul_20_sink_busy;
  wire _mul_20_busy;
  reg _mul_20_busy_reg;
  wire _mul_20_is_root;
  reg _mul_20_x_idle;
  reg [33-1:0] _mul_20_x_source_count;
  reg [5-1:0] _mul_20_x_source_mode;
  reg [16-1:0] _mul_20_x_source_generator_id;
  reg [32-1:0] _mul_20_x_source_offset;
  reg [33-1:0] _mul_20_x_source_size;
  reg [32-1:0] _mul_20_x_source_stride;
  reg [32-1:0] _mul_20_x_source_offset_buf;
  reg [33-1:0] _mul_20_x_source_size_buf;
  reg [32-1:0] _mul_20_x_source_stride_buf;
  reg [8-1:0] _mul_20_x_source_sel;
  reg [32-1:0] _mul_20_x_source_ram_raddr;
  reg _mul_20_x_source_ram_renable;
  wire [16-1:0] _mul_20_x_source_ram_rdata;
  reg _mul_20_x_source_fifo_deq;
  wire [16-1:0] _mul_20_x_source_fifo_rdata;
  reg [16-1:0] _mul_20_x_source_empty_data;
  reg _mul_20_y_idle;
  reg [33-1:0] _mul_20_y_source_count;
  reg [5-1:0] _mul_20_y_source_mode;
  reg [16-1:0] _mul_20_y_source_generator_id;
  reg [32-1:0] _mul_20_y_source_offset;
  reg [33-1:0] _mul_20_y_source_size;
  reg [32-1:0] _mul_20_y_source_stride;
  reg [32-1:0] _mul_20_y_source_offset_buf;
  reg [33-1:0] _mul_20_y_source_size_buf;
  reg [32-1:0] _mul_20_y_source_stride_buf;
  reg [8-1:0] _mul_20_y_source_sel;
  reg [32-1:0] _mul_20_y_source_ram_raddr;
  reg _mul_20_y_source_ram_renable;
  wire [16-1:0] _mul_20_y_source_ram_rdata;
  reg _mul_20_y_source_fifo_deq;
  wire [16-1:0] _mul_20_y_source_fifo_rdata;
  reg [16-1:0] _mul_20_y_source_empty_data;
  reg _mul_20_rshift_idle;
  reg [33-1:0] _mul_20_rshift_source_count;
  reg [5-1:0] _mul_20_rshift_source_mode;
  reg [16-1:0] _mul_20_rshift_source_generator_id;
  reg [32-1:0] _mul_20_rshift_source_offset;
  reg [33-1:0] _mul_20_rshift_source_size;
  reg [32-1:0] _mul_20_rshift_source_stride;
  reg [32-1:0] _mul_20_rshift_source_offset_buf;
  reg [33-1:0] _mul_20_rshift_source_size_buf;
  reg [32-1:0] _mul_20_rshift_source_stride_buf;
  reg [8-1:0] _mul_20_rshift_source_sel;
  reg [32-1:0] _mul_20_rshift_source_ram_raddr;
  reg _mul_20_rshift_source_ram_renable;
  wire [32-1:0] _mul_20_rshift_source_ram_rdata;
  reg _mul_20_rshift_source_fifo_deq;
  wire [32-1:0] _mul_20_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_20_rshift_source_empty_data;
  reg [33-1:0] _mul_20_z_sink_count;
  reg [5-1:0] _mul_20_z_sink_mode;
  reg [16-1:0] _mul_20_z_sink_generator_id;
  reg [32-1:0] _mul_20_z_sink_offset;
  reg [33-1:0] _mul_20_z_sink_size;
  reg [32-1:0] _mul_20_z_sink_stride;
  reg [32-1:0] _mul_20_z_sink_offset_buf;
  reg [33-1:0] _mul_20_z_sink_size_buf;
  reg [32-1:0] _mul_20_z_sink_stride_buf;
  reg [8-1:0] _mul_20_z_sink_sel;
  reg [32-1:0] _mul_20_z_sink_waddr;
  reg _mul_20_z_sink_wenable;
  reg [32-1:0] _mul_20_z_sink_wdata;
  reg _mul_20_z_sink_fifo_enq;
  reg [32-1:0] _mul_20_z_sink_fifo_wdata;
  reg [32-1:0] _mul_20_z_sink_immediate;
  reg _mul_21_stream_ivalid;
  wire _mul_21_stream_oready;
  wire _mul_21_stream_internal_oready;
  assign _mul_21_stream_internal_oready = 1;
  reg [32-1:0] _mul_21_fsm;
  localparam _mul_21_fsm_init = 0;
  wire _mul_21_run_flag;
  assign _mul_21_run_flag = 0;
  reg _mul_21_source_start;
  wire _mul_21_source_stop;
  reg _mul_21_source_busy;
  wire _mul_21_sink_start;
  wire _mul_21_sink_stop;
  wire _mul_21_sink_busy;
  wire _mul_21_busy;
  reg _mul_21_busy_reg;
  wire _mul_21_is_root;
  reg _mul_21_x_idle;
  reg [33-1:0] _mul_21_x_source_count;
  reg [5-1:0] _mul_21_x_source_mode;
  reg [16-1:0] _mul_21_x_source_generator_id;
  reg [32-1:0] _mul_21_x_source_offset;
  reg [33-1:0] _mul_21_x_source_size;
  reg [32-1:0] _mul_21_x_source_stride;
  reg [32-1:0] _mul_21_x_source_offset_buf;
  reg [33-1:0] _mul_21_x_source_size_buf;
  reg [32-1:0] _mul_21_x_source_stride_buf;
  reg [8-1:0] _mul_21_x_source_sel;
  reg [32-1:0] _mul_21_x_source_ram_raddr;
  reg _mul_21_x_source_ram_renable;
  wire [16-1:0] _mul_21_x_source_ram_rdata;
  reg _mul_21_x_source_fifo_deq;
  wire [16-1:0] _mul_21_x_source_fifo_rdata;
  reg [16-1:0] _mul_21_x_source_empty_data;
  reg _mul_21_y_idle;
  reg [33-1:0] _mul_21_y_source_count;
  reg [5-1:0] _mul_21_y_source_mode;
  reg [16-1:0] _mul_21_y_source_generator_id;
  reg [32-1:0] _mul_21_y_source_offset;
  reg [33-1:0] _mul_21_y_source_size;
  reg [32-1:0] _mul_21_y_source_stride;
  reg [32-1:0] _mul_21_y_source_offset_buf;
  reg [33-1:0] _mul_21_y_source_size_buf;
  reg [32-1:0] _mul_21_y_source_stride_buf;
  reg [8-1:0] _mul_21_y_source_sel;
  reg [32-1:0] _mul_21_y_source_ram_raddr;
  reg _mul_21_y_source_ram_renable;
  wire [16-1:0] _mul_21_y_source_ram_rdata;
  reg _mul_21_y_source_fifo_deq;
  wire [16-1:0] _mul_21_y_source_fifo_rdata;
  reg [16-1:0] _mul_21_y_source_empty_data;
  reg _mul_21_rshift_idle;
  reg [33-1:0] _mul_21_rshift_source_count;
  reg [5-1:0] _mul_21_rshift_source_mode;
  reg [16-1:0] _mul_21_rshift_source_generator_id;
  reg [32-1:0] _mul_21_rshift_source_offset;
  reg [33-1:0] _mul_21_rshift_source_size;
  reg [32-1:0] _mul_21_rshift_source_stride;
  reg [32-1:0] _mul_21_rshift_source_offset_buf;
  reg [33-1:0] _mul_21_rshift_source_size_buf;
  reg [32-1:0] _mul_21_rshift_source_stride_buf;
  reg [8-1:0] _mul_21_rshift_source_sel;
  reg [32-1:0] _mul_21_rshift_source_ram_raddr;
  reg _mul_21_rshift_source_ram_renable;
  wire [32-1:0] _mul_21_rshift_source_ram_rdata;
  reg _mul_21_rshift_source_fifo_deq;
  wire [32-1:0] _mul_21_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_21_rshift_source_empty_data;
  reg [33-1:0] _mul_21_z_sink_count;
  reg [5-1:0] _mul_21_z_sink_mode;
  reg [16-1:0] _mul_21_z_sink_generator_id;
  reg [32-1:0] _mul_21_z_sink_offset;
  reg [33-1:0] _mul_21_z_sink_size;
  reg [32-1:0] _mul_21_z_sink_stride;
  reg [32-1:0] _mul_21_z_sink_offset_buf;
  reg [33-1:0] _mul_21_z_sink_size_buf;
  reg [32-1:0] _mul_21_z_sink_stride_buf;
  reg [8-1:0] _mul_21_z_sink_sel;
  reg [32-1:0] _mul_21_z_sink_waddr;
  reg _mul_21_z_sink_wenable;
  reg [32-1:0] _mul_21_z_sink_wdata;
  reg _mul_21_z_sink_fifo_enq;
  reg [32-1:0] _mul_21_z_sink_fifo_wdata;
  reg [32-1:0] _mul_21_z_sink_immediate;
  reg _mul_22_stream_ivalid;
  wire _mul_22_stream_oready;
  wire _mul_22_stream_internal_oready;
  assign _mul_22_stream_internal_oready = 1;
  reg [32-1:0] _mul_22_fsm;
  localparam _mul_22_fsm_init = 0;
  wire _mul_22_run_flag;
  assign _mul_22_run_flag = 0;
  reg _mul_22_source_start;
  wire _mul_22_source_stop;
  reg _mul_22_source_busy;
  wire _mul_22_sink_start;
  wire _mul_22_sink_stop;
  wire _mul_22_sink_busy;
  wire _mul_22_busy;
  reg _mul_22_busy_reg;
  wire _mul_22_is_root;
  reg _mul_22_x_idle;
  reg [33-1:0] _mul_22_x_source_count;
  reg [5-1:0] _mul_22_x_source_mode;
  reg [16-1:0] _mul_22_x_source_generator_id;
  reg [32-1:0] _mul_22_x_source_offset;
  reg [33-1:0] _mul_22_x_source_size;
  reg [32-1:0] _mul_22_x_source_stride;
  reg [32-1:0] _mul_22_x_source_offset_buf;
  reg [33-1:0] _mul_22_x_source_size_buf;
  reg [32-1:0] _mul_22_x_source_stride_buf;
  reg [8-1:0] _mul_22_x_source_sel;
  reg [32-1:0] _mul_22_x_source_ram_raddr;
  reg _mul_22_x_source_ram_renable;
  wire [16-1:0] _mul_22_x_source_ram_rdata;
  reg _mul_22_x_source_fifo_deq;
  wire [16-1:0] _mul_22_x_source_fifo_rdata;
  reg [16-1:0] _mul_22_x_source_empty_data;
  reg _mul_22_y_idle;
  reg [33-1:0] _mul_22_y_source_count;
  reg [5-1:0] _mul_22_y_source_mode;
  reg [16-1:0] _mul_22_y_source_generator_id;
  reg [32-1:0] _mul_22_y_source_offset;
  reg [33-1:0] _mul_22_y_source_size;
  reg [32-1:0] _mul_22_y_source_stride;
  reg [32-1:0] _mul_22_y_source_offset_buf;
  reg [33-1:0] _mul_22_y_source_size_buf;
  reg [32-1:0] _mul_22_y_source_stride_buf;
  reg [8-1:0] _mul_22_y_source_sel;
  reg [32-1:0] _mul_22_y_source_ram_raddr;
  reg _mul_22_y_source_ram_renable;
  wire [16-1:0] _mul_22_y_source_ram_rdata;
  reg _mul_22_y_source_fifo_deq;
  wire [16-1:0] _mul_22_y_source_fifo_rdata;
  reg [16-1:0] _mul_22_y_source_empty_data;
  reg _mul_22_rshift_idle;
  reg [33-1:0] _mul_22_rshift_source_count;
  reg [5-1:0] _mul_22_rshift_source_mode;
  reg [16-1:0] _mul_22_rshift_source_generator_id;
  reg [32-1:0] _mul_22_rshift_source_offset;
  reg [33-1:0] _mul_22_rshift_source_size;
  reg [32-1:0] _mul_22_rshift_source_stride;
  reg [32-1:0] _mul_22_rshift_source_offset_buf;
  reg [33-1:0] _mul_22_rshift_source_size_buf;
  reg [32-1:0] _mul_22_rshift_source_stride_buf;
  reg [8-1:0] _mul_22_rshift_source_sel;
  reg [32-1:0] _mul_22_rshift_source_ram_raddr;
  reg _mul_22_rshift_source_ram_renable;
  wire [32-1:0] _mul_22_rshift_source_ram_rdata;
  reg _mul_22_rshift_source_fifo_deq;
  wire [32-1:0] _mul_22_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_22_rshift_source_empty_data;
  reg [33-1:0] _mul_22_z_sink_count;
  reg [5-1:0] _mul_22_z_sink_mode;
  reg [16-1:0] _mul_22_z_sink_generator_id;
  reg [32-1:0] _mul_22_z_sink_offset;
  reg [33-1:0] _mul_22_z_sink_size;
  reg [32-1:0] _mul_22_z_sink_stride;
  reg [32-1:0] _mul_22_z_sink_offset_buf;
  reg [33-1:0] _mul_22_z_sink_size_buf;
  reg [32-1:0] _mul_22_z_sink_stride_buf;
  reg [8-1:0] _mul_22_z_sink_sel;
  reg [32-1:0] _mul_22_z_sink_waddr;
  reg _mul_22_z_sink_wenable;
  reg [32-1:0] _mul_22_z_sink_wdata;
  reg _mul_22_z_sink_fifo_enq;
  reg [32-1:0] _mul_22_z_sink_fifo_wdata;
  reg [32-1:0] _mul_22_z_sink_immediate;
  reg _mul_23_stream_ivalid;
  wire _mul_23_stream_oready;
  wire _mul_23_stream_internal_oready;
  assign _mul_23_stream_internal_oready = 1;
  reg [32-1:0] _mul_23_fsm;
  localparam _mul_23_fsm_init = 0;
  wire _mul_23_run_flag;
  assign _mul_23_run_flag = 0;
  reg _mul_23_source_start;
  wire _mul_23_source_stop;
  reg _mul_23_source_busy;
  wire _mul_23_sink_start;
  wire _mul_23_sink_stop;
  wire _mul_23_sink_busy;
  wire _mul_23_busy;
  reg _mul_23_busy_reg;
  wire _mul_23_is_root;
  reg _mul_23_x_idle;
  reg [33-1:0] _mul_23_x_source_count;
  reg [5-1:0] _mul_23_x_source_mode;
  reg [16-1:0] _mul_23_x_source_generator_id;
  reg [32-1:0] _mul_23_x_source_offset;
  reg [33-1:0] _mul_23_x_source_size;
  reg [32-1:0] _mul_23_x_source_stride;
  reg [32-1:0] _mul_23_x_source_offset_buf;
  reg [33-1:0] _mul_23_x_source_size_buf;
  reg [32-1:0] _mul_23_x_source_stride_buf;
  reg [8-1:0] _mul_23_x_source_sel;
  reg [32-1:0] _mul_23_x_source_ram_raddr;
  reg _mul_23_x_source_ram_renable;
  wire [16-1:0] _mul_23_x_source_ram_rdata;
  reg _mul_23_x_source_fifo_deq;
  wire [16-1:0] _mul_23_x_source_fifo_rdata;
  reg [16-1:0] _mul_23_x_source_empty_data;
  reg _mul_23_y_idle;
  reg [33-1:0] _mul_23_y_source_count;
  reg [5-1:0] _mul_23_y_source_mode;
  reg [16-1:0] _mul_23_y_source_generator_id;
  reg [32-1:0] _mul_23_y_source_offset;
  reg [33-1:0] _mul_23_y_source_size;
  reg [32-1:0] _mul_23_y_source_stride;
  reg [32-1:0] _mul_23_y_source_offset_buf;
  reg [33-1:0] _mul_23_y_source_size_buf;
  reg [32-1:0] _mul_23_y_source_stride_buf;
  reg [8-1:0] _mul_23_y_source_sel;
  reg [32-1:0] _mul_23_y_source_ram_raddr;
  reg _mul_23_y_source_ram_renable;
  wire [16-1:0] _mul_23_y_source_ram_rdata;
  reg _mul_23_y_source_fifo_deq;
  wire [16-1:0] _mul_23_y_source_fifo_rdata;
  reg [16-1:0] _mul_23_y_source_empty_data;
  reg _mul_23_rshift_idle;
  reg [33-1:0] _mul_23_rshift_source_count;
  reg [5-1:0] _mul_23_rshift_source_mode;
  reg [16-1:0] _mul_23_rshift_source_generator_id;
  reg [32-1:0] _mul_23_rshift_source_offset;
  reg [33-1:0] _mul_23_rshift_source_size;
  reg [32-1:0] _mul_23_rshift_source_stride;
  reg [32-1:0] _mul_23_rshift_source_offset_buf;
  reg [33-1:0] _mul_23_rshift_source_size_buf;
  reg [32-1:0] _mul_23_rshift_source_stride_buf;
  reg [8-1:0] _mul_23_rshift_source_sel;
  reg [32-1:0] _mul_23_rshift_source_ram_raddr;
  reg _mul_23_rshift_source_ram_renable;
  wire [32-1:0] _mul_23_rshift_source_ram_rdata;
  reg _mul_23_rshift_source_fifo_deq;
  wire [32-1:0] _mul_23_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_23_rshift_source_empty_data;
  reg [33-1:0] _mul_23_z_sink_count;
  reg [5-1:0] _mul_23_z_sink_mode;
  reg [16-1:0] _mul_23_z_sink_generator_id;
  reg [32-1:0] _mul_23_z_sink_offset;
  reg [33-1:0] _mul_23_z_sink_size;
  reg [32-1:0] _mul_23_z_sink_stride;
  reg [32-1:0] _mul_23_z_sink_offset_buf;
  reg [33-1:0] _mul_23_z_sink_size_buf;
  reg [32-1:0] _mul_23_z_sink_stride_buf;
  reg [8-1:0] _mul_23_z_sink_sel;
  reg [32-1:0] _mul_23_z_sink_waddr;
  reg _mul_23_z_sink_wenable;
  reg [32-1:0] _mul_23_z_sink_wdata;
  reg _mul_23_z_sink_fifo_enq;
  reg [32-1:0] _mul_23_z_sink_fifo_wdata;
  reg [32-1:0] _mul_23_z_sink_immediate;
  reg _mul_24_stream_ivalid;
  wire _mul_24_stream_oready;
  wire _mul_24_stream_internal_oready;
  assign _mul_24_stream_internal_oready = 1;
  reg [32-1:0] _mul_24_fsm;
  localparam _mul_24_fsm_init = 0;
  wire _mul_24_run_flag;
  assign _mul_24_run_flag = 0;
  reg _mul_24_source_start;
  wire _mul_24_source_stop;
  reg _mul_24_source_busy;
  wire _mul_24_sink_start;
  wire _mul_24_sink_stop;
  wire _mul_24_sink_busy;
  wire _mul_24_busy;
  reg _mul_24_busy_reg;
  wire _mul_24_is_root;
  reg _mul_24_x_idle;
  reg [33-1:0] _mul_24_x_source_count;
  reg [5-1:0] _mul_24_x_source_mode;
  reg [16-1:0] _mul_24_x_source_generator_id;
  reg [32-1:0] _mul_24_x_source_offset;
  reg [33-1:0] _mul_24_x_source_size;
  reg [32-1:0] _mul_24_x_source_stride;
  reg [32-1:0] _mul_24_x_source_offset_buf;
  reg [33-1:0] _mul_24_x_source_size_buf;
  reg [32-1:0] _mul_24_x_source_stride_buf;
  reg [8-1:0] _mul_24_x_source_sel;
  reg [32-1:0] _mul_24_x_source_ram_raddr;
  reg _mul_24_x_source_ram_renable;
  wire [16-1:0] _mul_24_x_source_ram_rdata;
  reg _mul_24_x_source_fifo_deq;
  wire [16-1:0] _mul_24_x_source_fifo_rdata;
  reg [16-1:0] _mul_24_x_source_empty_data;
  reg _mul_24_y_idle;
  reg [33-1:0] _mul_24_y_source_count;
  reg [5-1:0] _mul_24_y_source_mode;
  reg [16-1:0] _mul_24_y_source_generator_id;
  reg [32-1:0] _mul_24_y_source_offset;
  reg [33-1:0] _mul_24_y_source_size;
  reg [32-1:0] _mul_24_y_source_stride;
  reg [32-1:0] _mul_24_y_source_offset_buf;
  reg [33-1:0] _mul_24_y_source_size_buf;
  reg [32-1:0] _mul_24_y_source_stride_buf;
  reg [8-1:0] _mul_24_y_source_sel;
  reg [32-1:0] _mul_24_y_source_ram_raddr;
  reg _mul_24_y_source_ram_renable;
  wire [16-1:0] _mul_24_y_source_ram_rdata;
  reg _mul_24_y_source_fifo_deq;
  wire [16-1:0] _mul_24_y_source_fifo_rdata;
  reg [16-1:0] _mul_24_y_source_empty_data;
  reg _mul_24_rshift_idle;
  reg [33-1:0] _mul_24_rshift_source_count;
  reg [5-1:0] _mul_24_rshift_source_mode;
  reg [16-1:0] _mul_24_rshift_source_generator_id;
  reg [32-1:0] _mul_24_rshift_source_offset;
  reg [33-1:0] _mul_24_rshift_source_size;
  reg [32-1:0] _mul_24_rshift_source_stride;
  reg [32-1:0] _mul_24_rshift_source_offset_buf;
  reg [33-1:0] _mul_24_rshift_source_size_buf;
  reg [32-1:0] _mul_24_rshift_source_stride_buf;
  reg [8-1:0] _mul_24_rshift_source_sel;
  reg [32-1:0] _mul_24_rshift_source_ram_raddr;
  reg _mul_24_rshift_source_ram_renable;
  wire [32-1:0] _mul_24_rshift_source_ram_rdata;
  reg _mul_24_rshift_source_fifo_deq;
  wire [32-1:0] _mul_24_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_24_rshift_source_empty_data;
  reg [33-1:0] _mul_24_z_sink_count;
  reg [5-1:0] _mul_24_z_sink_mode;
  reg [16-1:0] _mul_24_z_sink_generator_id;
  reg [32-1:0] _mul_24_z_sink_offset;
  reg [33-1:0] _mul_24_z_sink_size;
  reg [32-1:0] _mul_24_z_sink_stride;
  reg [32-1:0] _mul_24_z_sink_offset_buf;
  reg [33-1:0] _mul_24_z_sink_size_buf;
  reg [32-1:0] _mul_24_z_sink_stride_buf;
  reg [8-1:0] _mul_24_z_sink_sel;
  reg [32-1:0] _mul_24_z_sink_waddr;
  reg _mul_24_z_sink_wenable;
  reg [32-1:0] _mul_24_z_sink_wdata;
  reg _mul_24_z_sink_fifo_enq;
  reg [32-1:0] _mul_24_z_sink_fifo_wdata;
  reg [32-1:0] _mul_24_z_sink_immediate;
  reg _mul_25_stream_ivalid;
  wire _mul_25_stream_oready;
  wire _mul_25_stream_internal_oready;
  assign _mul_25_stream_internal_oready = 1;
  reg [32-1:0] _mul_25_fsm;
  localparam _mul_25_fsm_init = 0;
  wire _mul_25_run_flag;
  assign _mul_25_run_flag = 0;
  reg _mul_25_source_start;
  wire _mul_25_source_stop;
  reg _mul_25_source_busy;
  wire _mul_25_sink_start;
  wire _mul_25_sink_stop;
  wire _mul_25_sink_busy;
  wire _mul_25_busy;
  reg _mul_25_busy_reg;
  wire _mul_25_is_root;
  reg _mul_25_x_idle;
  reg [33-1:0] _mul_25_x_source_count;
  reg [5-1:0] _mul_25_x_source_mode;
  reg [16-1:0] _mul_25_x_source_generator_id;
  reg [32-1:0] _mul_25_x_source_offset;
  reg [33-1:0] _mul_25_x_source_size;
  reg [32-1:0] _mul_25_x_source_stride;
  reg [32-1:0] _mul_25_x_source_offset_buf;
  reg [33-1:0] _mul_25_x_source_size_buf;
  reg [32-1:0] _mul_25_x_source_stride_buf;
  reg [8-1:0] _mul_25_x_source_sel;
  reg [32-1:0] _mul_25_x_source_ram_raddr;
  reg _mul_25_x_source_ram_renable;
  wire [16-1:0] _mul_25_x_source_ram_rdata;
  reg _mul_25_x_source_fifo_deq;
  wire [16-1:0] _mul_25_x_source_fifo_rdata;
  reg [16-1:0] _mul_25_x_source_empty_data;
  reg _mul_25_y_idle;
  reg [33-1:0] _mul_25_y_source_count;
  reg [5-1:0] _mul_25_y_source_mode;
  reg [16-1:0] _mul_25_y_source_generator_id;
  reg [32-1:0] _mul_25_y_source_offset;
  reg [33-1:0] _mul_25_y_source_size;
  reg [32-1:0] _mul_25_y_source_stride;
  reg [32-1:0] _mul_25_y_source_offset_buf;
  reg [33-1:0] _mul_25_y_source_size_buf;
  reg [32-1:0] _mul_25_y_source_stride_buf;
  reg [8-1:0] _mul_25_y_source_sel;
  reg [32-1:0] _mul_25_y_source_ram_raddr;
  reg _mul_25_y_source_ram_renable;
  wire [16-1:0] _mul_25_y_source_ram_rdata;
  reg _mul_25_y_source_fifo_deq;
  wire [16-1:0] _mul_25_y_source_fifo_rdata;
  reg [16-1:0] _mul_25_y_source_empty_data;
  reg _mul_25_rshift_idle;
  reg [33-1:0] _mul_25_rshift_source_count;
  reg [5-1:0] _mul_25_rshift_source_mode;
  reg [16-1:0] _mul_25_rshift_source_generator_id;
  reg [32-1:0] _mul_25_rshift_source_offset;
  reg [33-1:0] _mul_25_rshift_source_size;
  reg [32-1:0] _mul_25_rshift_source_stride;
  reg [32-1:0] _mul_25_rshift_source_offset_buf;
  reg [33-1:0] _mul_25_rshift_source_size_buf;
  reg [32-1:0] _mul_25_rshift_source_stride_buf;
  reg [8-1:0] _mul_25_rshift_source_sel;
  reg [32-1:0] _mul_25_rshift_source_ram_raddr;
  reg _mul_25_rshift_source_ram_renable;
  wire [32-1:0] _mul_25_rshift_source_ram_rdata;
  reg _mul_25_rshift_source_fifo_deq;
  wire [32-1:0] _mul_25_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_25_rshift_source_empty_data;
  reg [33-1:0] _mul_25_z_sink_count;
  reg [5-1:0] _mul_25_z_sink_mode;
  reg [16-1:0] _mul_25_z_sink_generator_id;
  reg [32-1:0] _mul_25_z_sink_offset;
  reg [33-1:0] _mul_25_z_sink_size;
  reg [32-1:0] _mul_25_z_sink_stride;
  reg [32-1:0] _mul_25_z_sink_offset_buf;
  reg [33-1:0] _mul_25_z_sink_size_buf;
  reg [32-1:0] _mul_25_z_sink_stride_buf;
  reg [8-1:0] _mul_25_z_sink_sel;
  reg [32-1:0] _mul_25_z_sink_waddr;
  reg _mul_25_z_sink_wenable;
  reg [32-1:0] _mul_25_z_sink_wdata;
  reg _mul_25_z_sink_fifo_enq;
  reg [32-1:0] _mul_25_z_sink_fifo_wdata;
  reg [32-1:0] _mul_25_z_sink_immediate;
  reg _mul_26_stream_ivalid;
  wire _mul_26_stream_oready;
  wire _mul_26_stream_internal_oready;
  assign _mul_26_stream_internal_oready = 1;
  reg [32-1:0] _mul_26_fsm;
  localparam _mul_26_fsm_init = 0;
  wire _mul_26_run_flag;
  assign _mul_26_run_flag = 0;
  reg _mul_26_source_start;
  wire _mul_26_source_stop;
  reg _mul_26_source_busy;
  wire _mul_26_sink_start;
  wire _mul_26_sink_stop;
  wire _mul_26_sink_busy;
  wire _mul_26_busy;
  reg _mul_26_busy_reg;
  wire _mul_26_is_root;
  reg _mul_26_x_idle;
  reg [33-1:0] _mul_26_x_source_count;
  reg [5-1:0] _mul_26_x_source_mode;
  reg [16-1:0] _mul_26_x_source_generator_id;
  reg [32-1:0] _mul_26_x_source_offset;
  reg [33-1:0] _mul_26_x_source_size;
  reg [32-1:0] _mul_26_x_source_stride;
  reg [32-1:0] _mul_26_x_source_offset_buf;
  reg [33-1:0] _mul_26_x_source_size_buf;
  reg [32-1:0] _mul_26_x_source_stride_buf;
  reg [8-1:0] _mul_26_x_source_sel;
  reg [32-1:0] _mul_26_x_source_ram_raddr;
  reg _mul_26_x_source_ram_renable;
  wire [16-1:0] _mul_26_x_source_ram_rdata;
  reg _mul_26_x_source_fifo_deq;
  wire [16-1:0] _mul_26_x_source_fifo_rdata;
  reg [16-1:0] _mul_26_x_source_empty_data;
  reg _mul_26_y_idle;
  reg [33-1:0] _mul_26_y_source_count;
  reg [5-1:0] _mul_26_y_source_mode;
  reg [16-1:0] _mul_26_y_source_generator_id;
  reg [32-1:0] _mul_26_y_source_offset;
  reg [33-1:0] _mul_26_y_source_size;
  reg [32-1:0] _mul_26_y_source_stride;
  reg [32-1:0] _mul_26_y_source_offset_buf;
  reg [33-1:0] _mul_26_y_source_size_buf;
  reg [32-1:0] _mul_26_y_source_stride_buf;
  reg [8-1:0] _mul_26_y_source_sel;
  reg [32-1:0] _mul_26_y_source_ram_raddr;
  reg _mul_26_y_source_ram_renable;
  wire [16-1:0] _mul_26_y_source_ram_rdata;
  reg _mul_26_y_source_fifo_deq;
  wire [16-1:0] _mul_26_y_source_fifo_rdata;
  reg [16-1:0] _mul_26_y_source_empty_data;
  reg _mul_26_rshift_idle;
  reg [33-1:0] _mul_26_rshift_source_count;
  reg [5-1:0] _mul_26_rshift_source_mode;
  reg [16-1:0] _mul_26_rshift_source_generator_id;
  reg [32-1:0] _mul_26_rshift_source_offset;
  reg [33-1:0] _mul_26_rshift_source_size;
  reg [32-1:0] _mul_26_rshift_source_stride;
  reg [32-1:0] _mul_26_rshift_source_offset_buf;
  reg [33-1:0] _mul_26_rshift_source_size_buf;
  reg [32-1:0] _mul_26_rshift_source_stride_buf;
  reg [8-1:0] _mul_26_rshift_source_sel;
  reg [32-1:0] _mul_26_rshift_source_ram_raddr;
  reg _mul_26_rshift_source_ram_renable;
  wire [32-1:0] _mul_26_rshift_source_ram_rdata;
  reg _mul_26_rshift_source_fifo_deq;
  wire [32-1:0] _mul_26_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_26_rshift_source_empty_data;
  reg [33-1:0] _mul_26_z_sink_count;
  reg [5-1:0] _mul_26_z_sink_mode;
  reg [16-1:0] _mul_26_z_sink_generator_id;
  reg [32-1:0] _mul_26_z_sink_offset;
  reg [33-1:0] _mul_26_z_sink_size;
  reg [32-1:0] _mul_26_z_sink_stride;
  reg [32-1:0] _mul_26_z_sink_offset_buf;
  reg [33-1:0] _mul_26_z_sink_size_buf;
  reg [32-1:0] _mul_26_z_sink_stride_buf;
  reg [8-1:0] _mul_26_z_sink_sel;
  reg [32-1:0] _mul_26_z_sink_waddr;
  reg _mul_26_z_sink_wenable;
  reg [32-1:0] _mul_26_z_sink_wdata;
  reg _mul_26_z_sink_fifo_enq;
  reg [32-1:0] _mul_26_z_sink_fifo_wdata;
  reg [32-1:0] _mul_26_z_sink_immediate;
  reg _mul_27_stream_ivalid;
  wire _mul_27_stream_oready;
  wire _mul_27_stream_internal_oready;
  assign _mul_27_stream_internal_oready = 1;
  reg [32-1:0] _mul_27_fsm;
  localparam _mul_27_fsm_init = 0;
  wire _mul_27_run_flag;
  assign _mul_27_run_flag = 0;
  reg _mul_27_source_start;
  wire _mul_27_source_stop;
  reg _mul_27_source_busy;
  wire _mul_27_sink_start;
  wire _mul_27_sink_stop;
  wire _mul_27_sink_busy;
  wire _mul_27_busy;
  reg _mul_27_busy_reg;
  wire _mul_27_is_root;
  reg _mul_27_x_idle;
  reg [33-1:0] _mul_27_x_source_count;
  reg [5-1:0] _mul_27_x_source_mode;
  reg [16-1:0] _mul_27_x_source_generator_id;
  reg [32-1:0] _mul_27_x_source_offset;
  reg [33-1:0] _mul_27_x_source_size;
  reg [32-1:0] _mul_27_x_source_stride;
  reg [32-1:0] _mul_27_x_source_offset_buf;
  reg [33-1:0] _mul_27_x_source_size_buf;
  reg [32-1:0] _mul_27_x_source_stride_buf;
  reg [8-1:0] _mul_27_x_source_sel;
  reg [32-1:0] _mul_27_x_source_ram_raddr;
  reg _mul_27_x_source_ram_renable;
  wire [16-1:0] _mul_27_x_source_ram_rdata;
  reg _mul_27_x_source_fifo_deq;
  wire [16-1:0] _mul_27_x_source_fifo_rdata;
  reg [16-1:0] _mul_27_x_source_empty_data;
  reg _mul_27_y_idle;
  reg [33-1:0] _mul_27_y_source_count;
  reg [5-1:0] _mul_27_y_source_mode;
  reg [16-1:0] _mul_27_y_source_generator_id;
  reg [32-1:0] _mul_27_y_source_offset;
  reg [33-1:0] _mul_27_y_source_size;
  reg [32-1:0] _mul_27_y_source_stride;
  reg [32-1:0] _mul_27_y_source_offset_buf;
  reg [33-1:0] _mul_27_y_source_size_buf;
  reg [32-1:0] _mul_27_y_source_stride_buf;
  reg [8-1:0] _mul_27_y_source_sel;
  reg [32-1:0] _mul_27_y_source_ram_raddr;
  reg _mul_27_y_source_ram_renable;
  wire [16-1:0] _mul_27_y_source_ram_rdata;
  reg _mul_27_y_source_fifo_deq;
  wire [16-1:0] _mul_27_y_source_fifo_rdata;
  reg [16-1:0] _mul_27_y_source_empty_data;
  reg _mul_27_rshift_idle;
  reg [33-1:0] _mul_27_rshift_source_count;
  reg [5-1:0] _mul_27_rshift_source_mode;
  reg [16-1:0] _mul_27_rshift_source_generator_id;
  reg [32-1:0] _mul_27_rshift_source_offset;
  reg [33-1:0] _mul_27_rshift_source_size;
  reg [32-1:0] _mul_27_rshift_source_stride;
  reg [32-1:0] _mul_27_rshift_source_offset_buf;
  reg [33-1:0] _mul_27_rshift_source_size_buf;
  reg [32-1:0] _mul_27_rshift_source_stride_buf;
  reg [8-1:0] _mul_27_rshift_source_sel;
  reg [32-1:0] _mul_27_rshift_source_ram_raddr;
  reg _mul_27_rshift_source_ram_renable;
  wire [32-1:0] _mul_27_rshift_source_ram_rdata;
  reg _mul_27_rshift_source_fifo_deq;
  wire [32-1:0] _mul_27_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_27_rshift_source_empty_data;
  reg [33-1:0] _mul_27_z_sink_count;
  reg [5-1:0] _mul_27_z_sink_mode;
  reg [16-1:0] _mul_27_z_sink_generator_id;
  reg [32-1:0] _mul_27_z_sink_offset;
  reg [33-1:0] _mul_27_z_sink_size;
  reg [32-1:0] _mul_27_z_sink_stride;
  reg [32-1:0] _mul_27_z_sink_offset_buf;
  reg [33-1:0] _mul_27_z_sink_size_buf;
  reg [32-1:0] _mul_27_z_sink_stride_buf;
  reg [8-1:0] _mul_27_z_sink_sel;
  reg [32-1:0] _mul_27_z_sink_waddr;
  reg _mul_27_z_sink_wenable;
  reg [32-1:0] _mul_27_z_sink_wdata;
  reg _mul_27_z_sink_fifo_enq;
  reg [32-1:0] _mul_27_z_sink_fifo_wdata;
  reg [32-1:0] _mul_27_z_sink_immediate;
  reg _mul_28_stream_ivalid;
  wire _mul_28_stream_oready;
  wire _mul_28_stream_internal_oready;
  assign _mul_28_stream_internal_oready = 1;
  reg [32-1:0] _mul_28_fsm;
  localparam _mul_28_fsm_init = 0;
  wire _mul_28_run_flag;
  assign _mul_28_run_flag = 0;
  reg _mul_28_source_start;
  wire _mul_28_source_stop;
  reg _mul_28_source_busy;
  wire _mul_28_sink_start;
  wire _mul_28_sink_stop;
  wire _mul_28_sink_busy;
  wire _mul_28_busy;
  reg _mul_28_busy_reg;
  wire _mul_28_is_root;
  reg _mul_28_x_idle;
  reg [33-1:0] _mul_28_x_source_count;
  reg [5-1:0] _mul_28_x_source_mode;
  reg [16-1:0] _mul_28_x_source_generator_id;
  reg [32-1:0] _mul_28_x_source_offset;
  reg [33-1:0] _mul_28_x_source_size;
  reg [32-1:0] _mul_28_x_source_stride;
  reg [32-1:0] _mul_28_x_source_offset_buf;
  reg [33-1:0] _mul_28_x_source_size_buf;
  reg [32-1:0] _mul_28_x_source_stride_buf;
  reg [8-1:0] _mul_28_x_source_sel;
  reg [32-1:0] _mul_28_x_source_ram_raddr;
  reg _mul_28_x_source_ram_renable;
  wire [16-1:0] _mul_28_x_source_ram_rdata;
  reg _mul_28_x_source_fifo_deq;
  wire [16-1:0] _mul_28_x_source_fifo_rdata;
  reg [16-1:0] _mul_28_x_source_empty_data;
  reg _mul_28_y_idle;
  reg [33-1:0] _mul_28_y_source_count;
  reg [5-1:0] _mul_28_y_source_mode;
  reg [16-1:0] _mul_28_y_source_generator_id;
  reg [32-1:0] _mul_28_y_source_offset;
  reg [33-1:0] _mul_28_y_source_size;
  reg [32-1:0] _mul_28_y_source_stride;
  reg [32-1:0] _mul_28_y_source_offset_buf;
  reg [33-1:0] _mul_28_y_source_size_buf;
  reg [32-1:0] _mul_28_y_source_stride_buf;
  reg [8-1:0] _mul_28_y_source_sel;
  reg [32-1:0] _mul_28_y_source_ram_raddr;
  reg _mul_28_y_source_ram_renable;
  wire [16-1:0] _mul_28_y_source_ram_rdata;
  reg _mul_28_y_source_fifo_deq;
  wire [16-1:0] _mul_28_y_source_fifo_rdata;
  reg [16-1:0] _mul_28_y_source_empty_data;
  reg _mul_28_rshift_idle;
  reg [33-1:0] _mul_28_rshift_source_count;
  reg [5-1:0] _mul_28_rshift_source_mode;
  reg [16-1:0] _mul_28_rshift_source_generator_id;
  reg [32-1:0] _mul_28_rshift_source_offset;
  reg [33-1:0] _mul_28_rshift_source_size;
  reg [32-1:0] _mul_28_rshift_source_stride;
  reg [32-1:0] _mul_28_rshift_source_offset_buf;
  reg [33-1:0] _mul_28_rshift_source_size_buf;
  reg [32-1:0] _mul_28_rshift_source_stride_buf;
  reg [8-1:0] _mul_28_rshift_source_sel;
  reg [32-1:0] _mul_28_rshift_source_ram_raddr;
  reg _mul_28_rshift_source_ram_renable;
  wire [32-1:0] _mul_28_rshift_source_ram_rdata;
  reg _mul_28_rshift_source_fifo_deq;
  wire [32-1:0] _mul_28_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_28_rshift_source_empty_data;
  reg [33-1:0] _mul_28_z_sink_count;
  reg [5-1:0] _mul_28_z_sink_mode;
  reg [16-1:0] _mul_28_z_sink_generator_id;
  reg [32-1:0] _mul_28_z_sink_offset;
  reg [33-1:0] _mul_28_z_sink_size;
  reg [32-1:0] _mul_28_z_sink_stride;
  reg [32-1:0] _mul_28_z_sink_offset_buf;
  reg [33-1:0] _mul_28_z_sink_size_buf;
  reg [32-1:0] _mul_28_z_sink_stride_buf;
  reg [8-1:0] _mul_28_z_sink_sel;
  reg [32-1:0] _mul_28_z_sink_waddr;
  reg _mul_28_z_sink_wenable;
  reg [32-1:0] _mul_28_z_sink_wdata;
  reg _mul_28_z_sink_fifo_enq;
  reg [32-1:0] _mul_28_z_sink_fifo_wdata;
  reg [32-1:0] _mul_28_z_sink_immediate;
  reg _mul_29_stream_ivalid;
  wire _mul_29_stream_oready;
  wire _mul_29_stream_internal_oready;
  assign _mul_29_stream_internal_oready = 1;
  reg [32-1:0] _mul_29_fsm;
  localparam _mul_29_fsm_init = 0;
  wire _mul_29_run_flag;
  assign _mul_29_run_flag = 0;
  reg _mul_29_source_start;
  wire _mul_29_source_stop;
  reg _mul_29_source_busy;
  wire _mul_29_sink_start;
  wire _mul_29_sink_stop;
  wire _mul_29_sink_busy;
  wire _mul_29_busy;
  reg _mul_29_busy_reg;
  wire _mul_29_is_root;
  reg _mul_29_x_idle;
  reg [33-1:0] _mul_29_x_source_count;
  reg [5-1:0] _mul_29_x_source_mode;
  reg [16-1:0] _mul_29_x_source_generator_id;
  reg [32-1:0] _mul_29_x_source_offset;
  reg [33-1:0] _mul_29_x_source_size;
  reg [32-1:0] _mul_29_x_source_stride;
  reg [32-1:0] _mul_29_x_source_offset_buf;
  reg [33-1:0] _mul_29_x_source_size_buf;
  reg [32-1:0] _mul_29_x_source_stride_buf;
  reg [8-1:0] _mul_29_x_source_sel;
  reg [32-1:0] _mul_29_x_source_ram_raddr;
  reg _mul_29_x_source_ram_renable;
  wire [16-1:0] _mul_29_x_source_ram_rdata;
  reg _mul_29_x_source_fifo_deq;
  wire [16-1:0] _mul_29_x_source_fifo_rdata;
  reg [16-1:0] _mul_29_x_source_empty_data;
  reg _mul_29_y_idle;
  reg [33-1:0] _mul_29_y_source_count;
  reg [5-1:0] _mul_29_y_source_mode;
  reg [16-1:0] _mul_29_y_source_generator_id;
  reg [32-1:0] _mul_29_y_source_offset;
  reg [33-1:0] _mul_29_y_source_size;
  reg [32-1:0] _mul_29_y_source_stride;
  reg [32-1:0] _mul_29_y_source_offset_buf;
  reg [33-1:0] _mul_29_y_source_size_buf;
  reg [32-1:0] _mul_29_y_source_stride_buf;
  reg [8-1:0] _mul_29_y_source_sel;
  reg [32-1:0] _mul_29_y_source_ram_raddr;
  reg _mul_29_y_source_ram_renable;
  wire [16-1:0] _mul_29_y_source_ram_rdata;
  reg _mul_29_y_source_fifo_deq;
  wire [16-1:0] _mul_29_y_source_fifo_rdata;
  reg [16-1:0] _mul_29_y_source_empty_data;
  reg _mul_29_rshift_idle;
  reg [33-1:0] _mul_29_rshift_source_count;
  reg [5-1:0] _mul_29_rshift_source_mode;
  reg [16-1:0] _mul_29_rshift_source_generator_id;
  reg [32-1:0] _mul_29_rshift_source_offset;
  reg [33-1:0] _mul_29_rshift_source_size;
  reg [32-1:0] _mul_29_rshift_source_stride;
  reg [32-1:0] _mul_29_rshift_source_offset_buf;
  reg [33-1:0] _mul_29_rshift_source_size_buf;
  reg [32-1:0] _mul_29_rshift_source_stride_buf;
  reg [8-1:0] _mul_29_rshift_source_sel;
  reg [32-1:0] _mul_29_rshift_source_ram_raddr;
  reg _mul_29_rshift_source_ram_renable;
  wire [32-1:0] _mul_29_rshift_source_ram_rdata;
  reg _mul_29_rshift_source_fifo_deq;
  wire [32-1:0] _mul_29_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_29_rshift_source_empty_data;
  reg [33-1:0] _mul_29_z_sink_count;
  reg [5-1:0] _mul_29_z_sink_mode;
  reg [16-1:0] _mul_29_z_sink_generator_id;
  reg [32-1:0] _mul_29_z_sink_offset;
  reg [33-1:0] _mul_29_z_sink_size;
  reg [32-1:0] _mul_29_z_sink_stride;
  reg [32-1:0] _mul_29_z_sink_offset_buf;
  reg [33-1:0] _mul_29_z_sink_size_buf;
  reg [32-1:0] _mul_29_z_sink_stride_buf;
  reg [8-1:0] _mul_29_z_sink_sel;
  reg [32-1:0] _mul_29_z_sink_waddr;
  reg _mul_29_z_sink_wenable;
  reg [32-1:0] _mul_29_z_sink_wdata;
  reg _mul_29_z_sink_fifo_enq;
  reg [32-1:0] _mul_29_z_sink_fifo_wdata;
  reg [32-1:0] _mul_29_z_sink_immediate;
  reg _mul_30_stream_ivalid;
  wire _mul_30_stream_oready;
  wire _mul_30_stream_internal_oready;
  assign _mul_30_stream_internal_oready = 1;
  reg [32-1:0] _mul_30_fsm;
  localparam _mul_30_fsm_init = 0;
  wire _mul_30_run_flag;
  assign _mul_30_run_flag = 0;
  reg _mul_30_source_start;
  wire _mul_30_source_stop;
  reg _mul_30_source_busy;
  wire _mul_30_sink_start;
  wire _mul_30_sink_stop;
  wire _mul_30_sink_busy;
  wire _mul_30_busy;
  reg _mul_30_busy_reg;
  wire _mul_30_is_root;
  reg _mul_30_x_idle;
  reg [33-1:0] _mul_30_x_source_count;
  reg [5-1:0] _mul_30_x_source_mode;
  reg [16-1:0] _mul_30_x_source_generator_id;
  reg [32-1:0] _mul_30_x_source_offset;
  reg [33-1:0] _mul_30_x_source_size;
  reg [32-1:0] _mul_30_x_source_stride;
  reg [32-1:0] _mul_30_x_source_offset_buf;
  reg [33-1:0] _mul_30_x_source_size_buf;
  reg [32-1:0] _mul_30_x_source_stride_buf;
  reg [8-1:0] _mul_30_x_source_sel;
  reg [32-1:0] _mul_30_x_source_ram_raddr;
  reg _mul_30_x_source_ram_renable;
  wire [16-1:0] _mul_30_x_source_ram_rdata;
  reg _mul_30_x_source_fifo_deq;
  wire [16-1:0] _mul_30_x_source_fifo_rdata;
  reg [16-1:0] _mul_30_x_source_empty_data;
  reg _mul_30_y_idle;
  reg [33-1:0] _mul_30_y_source_count;
  reg [5-1:0] _mul_30_y_source_mode;
  reg [16-1:0] _mul_30_y_source_generator_id;
  reg [32-1:0] _mul_30_y_source_offset;
  reg [33-1:0] _mul_30_y_source_size;
  reg [32-1:0] _mul_30_y_source_stride;
  reg [32-1:0] _mul_30_y_source_offset_buf;
  reg [33-1:0] _mul_30_y_source_size_buf;
  reg [32-1:0] _mul_30_y_source_stride_buf;
  reg [8-1:0] _mul_30_y_source_sel;
  reg [32-1:0] _mul_30_y_source_ram_raddr;
  reg _mul_30_y_source_ram_renable;
  wire [16-1:0] _mul_30_y_source_ram_rdata;
  reg _mul_30_y_source_fifo_deq;
  wire [16-1:0] _mul_30_y_source_fifo_rdata;
  reg [16-1:0] _mul_30_y_source_empty_data;
  reg _mul_30_rshift_idle;
  reg [33-1:0] _mul_30_rshift_source_count;
  reg [5-1:0] _mul_30_rshift_source_mode;
  reg [16-1:0] _mul_30_rshift_source_generator_id;
  reg [32-1:0] _mul_30_rshift_source_offset;
  reg [33-1:0] _mul_30_rshift_source_size;
  reg [32-1:0] _mul_30_rshift_source_stride;
  reg [32-1:0] _mul_30_rshift_source_offset_buf;
  reg [33-1:0] _mul_30_rshift_source_size_buf;
  reg [32-1:0] _mul_30_rshift_source_stride_buf;
  reg [8-1:0] _mul_30_rshift_source_sel;
  reg [32-1:0] _mul_30_rshift_source_ram_raddr;
  reg _mul_30_rshift_source_ram_renable;
  wire [32-1:0] _mul_30_rshift_source_ram_rdata;
  reg _mul_30_rshift_source_fifo_deq;
  wire [32-1:0] _mul_30_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_30_rshift_source_empty_data;
  reg [33-1:0] _mul_30_z_sink_count;
  reg [5-1:0] _mul_30_z_sink_mode;
  reg [16-1:0] _mul_30_z_sink_generator_id;
  reg [32-1:0] _mul_30_z_sink_offset;
  reg [33-1:0] _mul_30_z_sink_size;
  reg [32-1:0] _mul_30_z_sink_stride;
  reg [32-1:0] _mul_30_z_sink_offset_buf;
  reg [33-1:0] _mul_30_z_sink_size_buf;
  reg [32-1:0] _mul_30_z_sink_stride_buf;
  reg [8-1:0] _mul_30_z_sink_sel;
  reg [32-1:0] _mul_30_z_sink_waddr;
  reg _mul_30_z_sink_wenable;
  reg [32-1:0] _mul_30_z_sink_wdata;
  reg _mul_30_z_sink_fifo_enq;
  reg [32-1:0] _mul_30_z_sink_fifo_wdata;
  reg [32-1:0] _mul_30_z_sink_immediate;
  reg _mul_31_stream_ivalid;
  wire _mul_31_stream_oready;
  wire _mul_31_stream_internal_oready;
  assign _mul_31_stream_internal_oready = 1;
  reg [32-1:0] _mul_31_fsm;
  localparam _mul_31_fsm_init = 0;
  wire _mul_31_run_flag;
  assign _mul_31_run_flag = 0;
  reg _mul_31_source_start;
  wire _mul_31_source_stop;
  reg _mul_31_source_busy;
  wire _mul_31_sink_start;
  wire _mul_31_sink_stop;
  wire _mul_31_sink_busy;
  wire _mul_31_busy;
  reg _mul_31_busy_reg;
  wire _mul_31_is_root;
  reg _mul_31_x_idle;
  reg [33-1:0] _mul_31_x_source_count;
  reg [5-1:0] _mul_31_x_source_mode;
  reg [16-1:0] _mul_31_x_source_generator_id;
  reg [32-1:0] _mul_31_x_source_offset;
  reg [33-1:0] _mul_31_x_source_size;
  reg [32-1:0] _mul_31_x_source_stride;
  reg [32-1:0] _mul_31_x_source_offset_buf;
  reg [33-1:0] _mul_31_x_source_size_buf;
  reg [32-1:0] _mul_31_x_source_stride_buf;
  reg [8-1:0] _mul_31_x_source_sel;
  reg [32-1:0] _mul_31_x_source_ram_raddr;
  reg _mul_31_x_source_ram_renable;
  wire [16-1:0] _mul_31_x_source_ram_rdata;
  reg _mul_31_x_source_fifo_deq;
  wire [16-1:0] _mul_31_x_source_fifo_rdata;
  reg [16-1:0] _mul_31_x_source_empty_data;
  reg _mul_31_y_idle;
  reg [33-1:0] _mul_31_y_source_count;
  reg [5-1:0] _mul_31_y_source_mode;
  reg [16-1:0] _mul_31_y_source_generator_id;
  reg [32-1:0] _mul_31_y_source_offset;
  reg [33-1:0] _mul_31_y_source_size;
  reg [32-1:0] _mul_31_y_source_stride;
  reg [32-1:0] _mul_31_y_source_offset_buf;
  reg [33-1:0] _mul_31_y_source_size_buf;
  reg [32-1:0] _mul_31_y_source_stride_buf;
  reg [8-1:0] _mul_31_y_source_sel;
  reg [32-1:0] _mul_31_y_source_ram_raddr;
  reg _mul_31_y_source_ram_renable;
  wire [16-1:0] _mul_31_y_source_ram_rdata;
  reg _mul_31_y_source_fifo_deq;
  wire [16-1:0] _mul_31_y_source_fifo_rdata;
  reg [16-1:0] _mul_31_y_source_empty_data;
  reg _mul_31_rshift_idle;
  reg [33-1:0] _mul_31_rshift_source_count;
  reg [5-1:0] _mul_31_rshift_source_mode;
  reg [16-1:0] _mul_31_rshift_source_generator_id;
  reg [32-1:0] _mul_31_rshift_source_offset;
  reg [33-1:0] _mul_31_rshift_source_size;
  reg [32-1:0] _mul_31_rshift_source_stride;
  reg [32-1:0] _mul_31_rshift_source_offset_buf;
  reg [33-1:0] _mul_31_rshift_source_size_buf;
  reg [32-1:0] _mul_31_rshift_source_stride_buf;
  reg [8-1:0] _mul_31_rshift_source_sel;
  reg [32-1:0] _mul_31_rshift_source_ram_raddr;
  reg _mul_31_rshift_source_ram_renable;
  wire [32-1:0] _mul_31_rshift_source_ram_rdata;
  reg _mul_31_rshift_source_fifo_deq;
  wire [32-1:0] _mul_31_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_31_rshift_source_empty_data;
  reg [33-1:0] _mul_31_z_sink_count;
  reg [5-1:0] _mul_31_z_sink_mode;
  reg [16-1:0] _mul_31_z_sink_generator_id;
  reg [32-1:0] _mul_31_z_sink_offset;
  reg [33-1:0] _mul_31_z_sink_size;
  reg [32-1:0] _mul_31_z_sink_stride;
  reg [32-1:0] _mul_31_z_sink_offset_buf;
  reg [33-1:0] _mul_31_z_sink_size_buf;
  reg [32-1:0] _mul_31_z_sink_stride_buf;
  reg [8-1:0] _mul_31_z_sink_sel;
  reg [32-1:0] _mul_31_z_sink_waddr;
  reg _mul_31_z_sink_wenable;
  reg [32-1:0] _mul_31_z_sink_wdata;
  reg _mul_31_z_sink_fifo_enq;
  reg [32-1:0] _mul_31_z_sink_fifo_wdata;
  reg [32-1:0] _mul_31_z_sink_immediate;
  reg _mul_32_stream_ivalid;
  wire _mul_32_stream_oready;
  wire _mul_32_stream_internal_oready;
  assign _mul_32_stream_internal_oready = 1;
  reg [32-1:0] _mul_32_fsm;
  localparam _mul_32_fsm_init = 0;
  wire _mul_32_run_flag;
  assign _mul_32_run_flag = 0;
  reg _mul_32_source_start;
  wire _mul_32_source_stop;
  reg _mul_32_source_busy;
  wire _mul_32_sink_start;
  wire _mul_32_sink_stop;
  wire _mul_32_sink_busy;
  wire _mul_32_busy;
  reg _mul_32_busy_reg;
  wire _mul_32_is_root;
  reg _mul_32_x_idle;
  reg [33-1:0] _mul_32_x_source_count;
  reg [5-1:0] _mul_32_x_source_mode;
  reg [16-1:0] _mul_32_x_source_generator_id;
  reg [32-1:0] _mul_32_x_source_offset;
  reg [33-1:0] _mul_32_x_source_size;
  reg [32-1:0] _mul_32_x_source_stride;
  reg [32-1:0] _mul_32_x_source_offset_buf;
  reg [33-1:0] _mul_32_x_source_size_buf;
  reg [32-1:0] _mul_32_x_source_stride_buf;
  reg [8-1:0] _mul_32_x_source_sel;
  reg [32-1:0] _mul_32_x_source_ram_raddr;
  reg _mul_32_x_source_ram_renable;
  wire [16-1:0] _mul_32_x_source_ram_rdata;
  reg _mul_32_x_source_fifo_deq;
  wire [16-1:0] _mul_32_x_source_fifo_rdata;
  reg [16-1:0] _mul_32_x_source_empty_data;
  reg _mul_32_y_idle;
  reg [33-1:0] _mul_32_y_source_count;
  reg [5-1:0] _mul_32_y_source_mode;
  reg [16-1:0] _mul_32_y_source_generator_id;
  reg [32-1:0] _mul_32_y_source_offset;
  reg [33-1:0] _mul_32_y_source_size;
  reg [32-1:0] _mul_32_y_source_stride;
  reg [32-1:0] _mul_32_y_source_offset_buf;
  reg [33-1:0] _mul_32_y_source_size_buf;
  reg [32-1:0] _mul_32_y_source_stride_buf;
  reg [8-1:0] _mul_32_y_source_sel;
  reg [32-1:0] _mul_32_y_source_ram_raddr;
  reg _mul_32_y_source_ram_renable;
  wire [16-1:0] _mul_32_y_source_ram_rdata;
  reg _mul_32_y_source_fifo_deq;
  wire [16-1:0] _mul_32_y_source_fifo_rdata;
  reg [16-1:0] _mul_32_y_source_empty_data;
  reg _mul_32_rshift_idle;
  reg [33-1:0] _mul_32_rshift_source_count;
  reg [5-1:0] _mul_32_rshift_source_mode;
  reg [16-1:0] _mul_32_rshift_source_generator_id;
  reg [32-1:0] _mul_32_rshift_source_offset;
  reg [33-1:0] _mul_32_rshift_source_size;
  reg [32-1:0] _mul_32_rshift_source_stride;
  reg [32-1:0] _mul_32_rshift_source_offset_buf;
  reg [33-1:0] _mul_32_rshift_source_size_buf;
  reg [32-1:0] _mul_32_rshift_source_stride_buf;
  reg [8-1:0] _mul_32_rshift_source_sel;
  reg [32-1:0] _mul_32_rshift_source_ram_raddr;
  reg _mul_32_rshift_source_ram_renable;
  wire [32-1:0] _mul_32_rshift_source_ram_rdata;
  reg _mul_32_rshift_source_fifo_deq;
  wire [32-1:0] _mul_32_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_32_rshift_source_empty_data;
  reg [33-1:0] _mul_32_z_sink_count;
  reg [5-1:0] _mul_32_z_sink_mode;
  reg [16-1:0] _mul_32_z_sink_generator_id;
  reg [32-1:0] _mul_32_z_sink_offset;
  reg [33-1:0] _mul_32_z_sink_size;
  reg [32-1:0] _mul_32_z_sink_stride;
  reg [32-1:0] _mul_32_z_sink_offset_buf;
  reg [33-1:0] _mul_32_z_sink_size_buf;
  reg [32-1:0] _mul_32_z_sink_stride_buf;
  reg [8-1:0] _mul_32_z_sink_sel;
  reg [32-1:0] _mul_32_z_sink_waddr;
  reg _mul_32_z_sink_wenable;
  reg [32-1:0] _mul_32_z_sink_wdata;
  reg _mul_32_z_sink_fifo_enq;
  reg [32-1:0] _mul_32_z_sink_fifo_wdata;
  reg [32-1:0] _mul_32_z_sink_immediate;
  reg _mul_33_stream_ivalid;
  wire _mul_33_stream_oready;
  wire _mul_33_stream_internal_oready;
  assign _mul_33_stream_internal_oready = 1;
  reg [32-1:0] _mul_33_fsm;
  localparam _mul_33_fsm_init = 0;
  wire _mul_33_run_flag;
  assign _mul_33_run_flag = 0;
  reg _mul_33_source_start;
  wire _mul_33_source_stop;
  reg _mul_33_source_busy;
  wire _mul_33_sink_start;
  wire _mul_33_sink_stop;
  wire _mul_33_sink_busy;
  wire _mul_33_busy;
  reg _mul_33_busy_reg;
  wire _mul_33_is_root;
  reg _mul_33_x_idle;
  reg [33-1:0] _mul_33_x_source_count;
  reg [5-1:0] _mul_33_x_source_mode;
  reg [16-1:0] _mul_33_x_source_generator_id;
  reg [32-1:0] _mul_33_x_source_offset;
  reg [33-1:0] _mul_33_x_source_size;
  reg [32-1:0] _mul_33_x_source_stride;
  reg [32-1:0] _mul_33_x_source_offset_buf;
  reg [33-1:0] _mul_33_x_source_size_buf;
  reg [32-1:0] _mul_33_x_source_stride_buf;
  reg [8-1:0] _mul_33_x_source_sel;
  reg [32-1:0] _mul_33_x_source_ram_raddr;
  reg _mul_33_x_source_ram_renable;
  wire [16-1:0] _mul_33_x_source_ram_rdata;
  reg _mul_33_x_source_fifo_deq;
  wire [16-1:0] _mul_33_x_source_fifo_rdata;
  reg [16-1:0] _mul_33_x_source_empty_data;
  reg _mul_33_y_idle;
  reg [33-1:0] _mul_33_y_source_count;
  reg [5-1:0] _mul_33_y_source_mode;
  reg [16-1:0] _mul_33_y_source_generator_id;
  reg [32-1:0] _mul_33_y_source_offset;
  reg [33-1:0] _mul_33_y_source_size;
  reg [32-1:0] _mul_33_y_source_stride;
  reg [32-1:0] _mul_33_y_source_offset_buf;
  reg [33-1:0] _mul_33_y_source_size_buf;
  reg [32-1:0] _mul_33_y_source_stride_buf;
  reg [8-1:0] _mul_33_y_source_sel;
  reg [32-1:0] _mul_33_y_source_ram_raddr;
  reg _mul_33_y_source_ram_renable;
  wire [16-1:0] _mul_33_y_source_ram_rdata;
  reg _mul_33_y_source_fifo_deq;
  wire [16-1:0] _mul_33_y_source_fifo_rdata;
  reg [16-1:0] _mul_33_y_source_empty_data;
  reg _mul_33_rshift_idle;
  reg [33-1:0] _mul_33_rshift_source_count;
  reg [5-1:0] _mul_33_rshift_source_mode;
  reg [16-1:0] _mul_33_rshift_source_generator_id;
  reg [32-1:0] _mul_33_rshift_source_offset;
  reg [33-1:0] _mul_33_rshift_source_size;
  reg [32-1:0] _mul_33_rshift_source_stride;
  reg [32-1:0] _mul_33_rshift_source_offset_buf;
  reg [33-1:0] _mul_33_rshift_source_size_buf;
  reg [32-1:0] _mul_33_rshift_source_stride_buf;
  reg [8-1:0] _mul_33_rshift_source_sel;
  reg [32-1:0] _mul_33_rshift_source_ram_raddr;
  reg _mul_33_rshift_source_ram_renable;
  wire [32-1:0] _mul_33_rshift_source_ram_rdata;
  reg _mul_33_rshift_source_fifo_deq;
  wire [32-1:0] _mul_33_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_33_rshift_source_empty_data;
  reg [33-1:0] _mul_33_z_sink_count;
  reg [5-1:0] _mul_33_z_sink_mode;
  reg [16-1:0] _mul_33_z_sink_generator_id;
  reg [32-1:0] _mul_33_z_sink_offset;
  reg [33-1:0] _mul_33_z_sink_size;
  reg [32-1:0] _mul_33_z_sink_stride;
  reg [32-1:0] _mul_33_z_sink_offset_buf;
  reg [33-1:0] _mul_33_z_sink_size_buf;
  reg [32-1:0] _mul_33_z_sink_stride_buf;
  reg [8-1:0] _mul_33_z_sink_sel;
  reg [32-1:0] _mul_33_z_sink_waddr;
  reg _mul_33_z_sink_wenable;
  reg [32-1:0] _mul_33_z_sink_wdata;
  reg _mul_33_z_sink_fifo_enq;
  reg [32-1:0] _mul_33_z_sink_fifo_wdata;
  reg [32-1:0] _mul_33_z_sink_immediate;
  reg _mul_34_stream_ivalid;
  wire _mul_34_stream_oready;
  wire _mul_34_stream_internal_oready;
  assign _mul_34_stream_internal_oready = 1;
  reg [32-1:0] _mul_34_fsm;
  localparam _mul_34_fsm_init = 0;
  wire _mul_34_run_flag;
  assign _mul_34_run_flag = 0;
  reg _mul_34_source_start;
  wire _mul_34_source_stop;
  reg _mul_34_source_busy;
  wire _mul_34_sink_start;
  wire _mul_34_sink_stop;
  wire _mul_34_sink_busy;
  wire _mul_34_busy;
  reg _mul_34_busy_reg;
  wire _mul_34_is_root;
  reg _mul_34_x_idle;
  reg [33-1:0] _mul_34_x_source_count;
  reg [5-1:0] _mul_34_x_source_mode;
  reg [16-1:0] _mul_34_x_source_generator_id;
  reg [32-1:0] _mul_34_x_source_offset;
  reg [33-1:0] _mul_34_x_source_size;
  reg [32-1:0] _mul_34_x_source_stride;
  reg [32-1:0] _mul_34_x_source_offset_buf;
  reg [33-1:0] _mul_34_x_source_size_buf;
  reg [32-1:0] _mul_34_x_source_stride_buf;
  reg [8-1:0] _mul_34_x_source_sel;
  reg [32-1:0] _mul_34_x_source_ram_raddr;
  reg _mul_34_x_source_ram_renable;
  wire [16-1:0] _mul_34_x_source_ram_rdata;
  reg _mul_34_x_source_fifo_deq;
  wire [16-1:0] _mul_34_x_source_fifo_rdata;
  reg [16-1:0] _mul_34_x_source_empty_data;
  reg _mul_34_y_idle;
  reg [33-1:0] _mul_34_y_source_count;
  reg [5-1:0] _mul_34_y_source_mode;
  reg [16-1:0] _mul_34_y_source_generator_id;
  reg [32-1:0] _mul_34_y_source_offset;
  reg [33-1:0] _mul_34_y_source_size;
  reg [32-1:0] _mul_34_y_source_stride;
  reg [32-1:0] _mul_34_y_source_offset_buf;
  reg [33-1:0] _mul_34_y_source_size_buf;
  reg [32-1:0] _mul_34_y_source_stride_buf;
  reg [8-1:0] _mul_34_y_source_sel;
  reg [32-1:0] _mul_34_y_source_ram_raddr;
  reg _mul_34_y_source_ram_renable;
  wire [16-1:0] _mul_34_y_source_ram_rdata;
  reg _mul_34_y_source_fifo_deq;
  wire [16-1:0] _mul_34_y_source_fifo_rdata;
  reg [16-1:0] _mul_34_y_source_empty_data;
  reg _mul_34_rshift_idle;
  reg [33-1:0] _mul_34_rshift_source_count;
  reg [5-1:0] _mul_34_rshift_source_mode;
  reg [16-1:0] _mul_34_rshift_source_generator_id;
  reg [32-1:0] _mul_34_rshift_source_offset;
  reg [33-1:0] _mul_34_rshift_source_size;
  reg [32-1:0] _mul_34_rshift_source_stride;
  reg [32-1:0] _mul_34_rshift_source_offset_buf;
  reg [33-1:0] _mul_34_rshift_source_size_buf;
  reg [32-1:0] _mul_34_rshift_source_stride_buf;
  reg [8-1:0] _mul_34_rshift_source_sel;
  reg [32-1:0] _mul_34_rshift_source_ram_raddr;
  reg _mul_34_rshift_source_ram_renable;
  wire [32-1:0] _mul_34_rshift_source_ram_rdata;
  reg _mul_34_rshift_source_fifo_deq;
  wire [32-1:0] _mul_34_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_34_rshift_source_empty_data;
  reg [33-1:0] _mul_34_z_sink_count;
  reg [5-1:0] _mul_34_z_sink_mode;
  reg [16-1:0] _mul_34_z_sink_generator_id;
  reg [32-1:0] _mul_34_z_sink_offset;
  reg [33-1:0] _mul_34_z_sink_size;
  reg [32-1:0] _mul_34_z_sink_stride;
  reg [32-1:0] _mul_34_z_sink_offset_buf;
  reg [33-1:0] _mul_34_z_sink_size_buf;
  reg [32-1:0] _mul_34_z_sink_stride_buf;
  reg [8-1:0] _mul_34_z_sink_sel;
  reg [32-1:0] _mul_34_z_sink_waddr;
  reg _mul_34_z_sink_wenable;
  reg [32-1:0] _mul_34_z_sink_wdata;
  reg _mul_34_z_sink_fifo_enq;
  reg [32-1:0] _mul_34_z_sink_fifo_wdata;
  reg [32-1:0] _mul_34_z_sink_immediate;
  reg _mul_35_stream_ivalid;
  wire _mul_35_stream_oready;
  wire _mul_35_stream_internal_oready;
  assign _mul_35_stream_internal_oready = 1;
  reg [32-1:0] _mul_35_fsm;
  localparam _mul_35_fsm_init = 0;
  wire _mul_35_run_flag;
  assign _mul_35_run_flag = 0;
  reg _mul_35_source_start;
  wire _mul_35_source_stop;
  reg _mul_35_source_busy;
  wire _mul_35_sink_start;
  wire _mul_35_sink_stop;
  wire _mul_35_sink_busy;
  wire _mul_35_busy;
  reg _mul_35_busy_reg;
  wire _mul_35_is_root;
  reg _mul_35_x_idle;
  reg [33-1:0] _mul_35_x_source_count;
  reg [5-1:0] _mul_35_x_source_mode;
  reg [16-1:0] _mul_35_x_source_generator_id;
  reg [32-1:0] _mul_35_x_source_offset;
  reg [33-1:0] _mul_35_x_source_size;
  reg [32-1:0] _mul_35_x_source_stride;
  reg [32-1:0] _mul_35_x_source_offset_buf;
  reg [33-1:0] _mul_35_x_source_size_buf;
  reg [32-1:0] _mul_35_x_source_stride_buf;
  reg [8-1:0] _mul_35_x_source_sel;
  reg [32-1:0] _mul_35_x_source_ram_raddr;
  reg _mul_35_x_source_ram_renable;
  wire [16-1:0] _mul_35_x_source_ram_rdata;
  reg _mul_35_x_source_fifo_deq;
  wire [16-1:0] _mul_35_x_source_fifo_rdata;
  reg [16-1:0] _mul_35_x_source_empty_data;
  reg _mul_35_y_idle;
  reg [33-1:0] _mul_35_y_source_count;
  reg [5-1:0] _mul_35_y_source_mode;
  reg [16-1:0] _mul_35_y_source_generator_id;
  reg [32-1:0] _mul_35_y_source_offset;
  reg [33-1:0] _mul_35_y_source_size;
  reg [32-1:0] _mul_35_y_source_stride;
  reg [32-1:0] _mul_35_y_source_offset_buf;
  reg [33-1:0] _mul_35_y_source_size_buf;
  reg [32-1:0] _mul_35_y_source_stride_buf;
  reg [8-1:0] _mul_35_y_source_sel;
  reg [32-1:0] _mul_35_y_source_ram_raddr;
  reg _mul_35_y_source_ram_renable;
  wire [16-1:0] _mul_35_y_source_ram_rdata;
  reg _mul_35_y_source_fifo_deq;
  wire [16-1:0] _mul_35_y_source_fifo_rdata;
  reg [16-1:0] _mul_35_y_source_empty_data;
  reg _mul_35_rshift_idle;
  reg [33-1:0] _mul_35_rshift_source_count;
  reg [5-1:0] _mul_35_rshift_source_mode;
  reg [16-1:0] _mul_35_rshift_source_generator_id;
  reg [32-1:0] _mul_35_rshift_source_offset;
  reg [33-1:0] _mul_35_rshift_source_size;
  reg [32-1:0] _mul_35_rshift_source_stride;
  reg [32-1:0] _mul_35_rshift_source_offset_buf;
  reg [33-1:0] _mul_35_rshift_source_size_buf;
  reg [32-1:0] _mul_35_rshift_source_stride_buf;
  reg [8-1:0] _mul_35_rshift_source_sel;
  reg [32-1:0] _mul_35_rshift_source_ram_raddr;
  reg _mul_35_rshift_source_ram_renable;
  wire [32-1:0] _mul_35_rshift_source_ram_rdata;
  reg _mul_35_rshift_source_fifo_deq;
  wire [32-1:0] _mul_35_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_35_rshift_source_empty_data;
  reg [33-1:0] _mul_35_z_sink_count;
  reg [5-1:0] _mul_35_z_sink_mode;
  reg [16-1:0] _mul_35_z_sink_generator_id;
  reg [32-1:0] _mul_35_z_sink_offset;
  reg [33-1:0] _mul_35_z_sink_size;
  reg [32-1:0] _mul_35_z_sink_stride;
  reg [32-1:0] _mul_35_z_sink_offset_buf;
  reg [33-1:0] _mul_35_z_sink_size_buf;
  reg [32-1:0] _mul_35_z_sink_stride_buf;
  reg [8-1:0] _mul_35_z_sink_sel;
  reg [32-1:0] _mul_35_z_sink_waddr;
  reg _mul_35_z_sink_wenable;
  reg [32-1:0] _mul_35_z_sink_wdata;
  reg _mul_35_z_sink_fifo_enq;
  reg [32-1:0] _mul_35_z_sink_fifo_wdata;
  reg [32-1:0] _mul_35_z_sink_immediate;
  reg _mul_36_stream_ivalid;
  wire _mul_36_stream_oready;
  wire _mul_36_stream_internal_oready;
  assign _mul_36_stream_internal_oready = 1;
  reg [32-1:0] _mul_36_fsm;
  localparam _mul_36_fsm_init = 0;
  wire _mul_36_run_flag;
  assign _mul_36_run_flag = 0;
  reg _mul_36_source_start;
  wire _mul_36_source_stop;
  reg _mul_36_source_busy;
  wire _mul_36_sink_start;
  wire _mul_36_sink_stop;
  wire _mul_36_sink_busy;
  wire _mul_36_busy;
  reg _mul_36_busy_reg;
  wire _mul_36_is_root;
  reg _mul_36_x_idle;
  reg [33-1:0] _mul_36_x_source_count;
  reg [5-1:0] _mul_36_x_source_mode;
  reg [16-1:0] _mul_36_x_source_generator_id;
  reg [32-1:0] _mul_36_x_source_offset;
  reg [33-1:0] _mul_36_x_source_size;
  reg [32-1:0] _mul_36_x_source_stride;
  reg [32-1:0] _mul_36_x_source_offset_buf;
  reg [33-1:0] _mul_36_x_source_size_buf;
  reg [32-1:0] _mul_36_x_source_stride_buf;
  reg [8-1:0] _mul_36_x_source_sel;
  reg [32-1:0] _mul_36_x_source_ram_raddr;
  reg _mul_36_x_source_ram_renable;
  wire [16-1:0] _mul_36_x_source_ram_rdata;
  reg _mul_36_x_source_fifo_deq;
  wire [16-1:0] _mul_36_x_source_fifo_rdata;
  reg [16-1:0] _mul_36_x_source_empty_data;
  reg _mul_36_y_idle;
  reg [33-1:0] _mul_36_y_source_count;
  reg [5-1:0] _mul_36_y_source_mode;
  reg [16-1:0] _mul_36_y_source_generator_id;
  reg [32-1:0] _mul_36_y_source_offset;
  reg [33-1:0] _mul_36_y_source_size;
  reg [32-1:0] _mul_36_y_source_stride;
  reg [32-1:0] _mul_36_y_source_offset_buf;
  reg [33-1:0] _mul_36_y_source_size_buf;
  reg [32-1:0] _mul_36_y_source_stride_buf;
  reg [8-1:0] _mul_36_y_source_sel;
  reg [32-1:0] _mul_36_y_source_ram_raddr;
  reg _mul_36_y_source_ram_renable;
  wire [16-1:0] _mul_36_y_source_ram_rdata;
  reg _mul_36_y_source_fifo_deq;
  wire [16-1:0] _mul_36_y_source_fifo_rdata;
  reg [16-1:0] _mul_36_y_source_empty_data;
  reg _mul_36_rshift_idle;
  reg [33-1:0] _mul_36_rshift_source_count;
  reg [5-1:0] _mul_36_rshift_source_mode;
  reg [16-1:0] _mul_36_rshift_source_generator_id;
  reg [32-1:0] _mul_36_rshift_source_offset;
  reg [33-1:0] _mul_36_rshift_source_size;
  reg [32-1:0] _mul_36_rshift_source_stride;
  reg [32-1:0] _mul_36_rshift_source_offset_buf;
  reg [33-1:0] _mul_36_rshift_source_size_buf;
  reg [32-1:0] _mul_36_rshift_source_stride_buf;
  reg [8-1:0] _mul_36_rshift_source_sel;
  reg [32-1:0] _mul_36_rshift_source_ram_raddr;
  reg _mul_36_rshift_source_ram_renable;
  wire [32-1:0] _mul_36_rshift_source_ram_rdata;
  reg _mul_36_rshift_source_fifo_deq;
  wire [32-1:0] _mul_36_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_36_rshift_source_empty_data;
  reg [33-1:0] _mul_36_z_sink_count;
  reg [5-1:0] _mul_36_z_sink_mode;
  reg [16-1:0] _mul_36_z_sink_generator_id;
  reg [32-1:0] _mul_36_z_sink_offset;
  reg [33-1:0] _mul_36_z_sink_size;
  reg [32-1:0] _mul_36_z_sink_stride;
  reg [32-1:0] _mul_36_z_sink_offset_buf;
  reg [33-1:0] _mul_36_z_sink_size_buf;
  reg [32-1:0] _mul_36_z_sink_stride_buf;
  reg [8-1:0] _mul_36_z_sink_sel;
  reg [32-1:0] _mul_36_z_sink_waddr;
  reg _mul_36_z_sink_wenable;
  reg [32-1:0] _mul_36_z_sink_wdata;
  reg _mul_36_z_sink_fifo_enq;
  reg [32-1:0] _mul_36_z_sink_fifo_wdata;
  reg [32-1:0] _mul_36_z_sink_immediate;
  reg _mul_37_stream_ivalid;
  wire _mul_37_stream_oready;
  wire _mul_37_stream_internal_oready;
  assign _mul_37_stream_internal_oready = 1;
  reg [32-1:0] _mul_37_fsm;
  localparam _mul_37_fsm_init = 0;
  wire _mul_37_run_flag;
  assign _mul_37_run_flag = 0;
  reg _mul_37_source_start;
  wire _mul_37_source_stop;
  reg _mul_37_source_busy;
  wire _mul_37_sink_start;
  wire _mul_37_sink_stop;
  wire _mul_37_sink_busy;
  wire _mul_37_busy;
  reg _mul_37_busy_reg;
  wire _mul_37_is_root;
  reg _mul_37_x_idle;
  reg [33-1:0] _mul_37_x_source_count;
  reg [5-1:0] _mul_37_x_source_mode;
  reg [16-1:0] _mul_37_x_source_generator_id;
  reg [32-1:0] _mul_37_x_source_offset;
  reg [33-1:0] _mul_37_x_source_size;
  reg [32-1:0] _mul_37_x_source_stride;
  reg [32-1:0] _mul_37_x_source_offset_buf;
  reg [33-1:0] _mul_37_x_source_size_buf;
  reg [32-1:0] _mul_37_x_source_stride_buf;
  reg [8-1:0] _mul_37_x_source_sel;
  reg [32-1:0] _mul_37_x_source_ram_raddr;
  reg _mul_37_x_source_ram_renable;
  wire [16-1:0] _mul_37_x_source_ram_rdata;
  reg _mul_37_x_source_fifo_deq;
  wire [16-1:0] _mul_37_x_source_fifo_rdata;
  reg [16-1:0] _mul_37_x_source_empty_data;
  reg _mul_37_y_idle;
  reg [33-1:0] _mul_37_y_source_count;
  reg [5-1:0] _mul_37_y_source_mode;
  reg [16-1:0] _mul_37_y_source_generator_id;
  reg [32-1:0] _mul_37_y_source_offset;
  reg [33-1:0] _mul_37_y_source_size;
  reg [32-1:0] _mul_37_y_source_stride;
  reg [32-1:0] _mul_37_y_source_offset_buf;
  reg [33-1:0] _mul_37_y_source_size_buf;
  reg [32-1:0] _mul_37_y_source_stride_buf;
  reg [8-1:0] _mul_37_y_source_sel;
  reg [32-1:0] _mul_37_y_source_ram_raddr;
  reg _mul_37_y_source_ram_renable;
  wire [16-1:0] _mul_37_y_source_ram_rdata;
  reg _mul_37_y_source_fifo_deq;
  wire [16-1:0] _mul_37_y_source_fifo_rdata;
  reg [16-1:0] _mul_37_y_source_empty_data;
  reg _mul_37_rshift_idle;
  reg [33-1:0] _mul_37_rshift_source_count;
  reg [5-1:0] _mul_37_rshift_source_mode;
  reg [16-1:0] _mul_37_rshift_source_generator_id;
  reg [32-1:0] _mul_37_rshift_source_offset;
  reg [33-1:0] _mul_37_rshift_source_size;
  reg [32-1:0] _mul_37_rshift_source_stride;
  reg [32-1:0] _mul_37_rshift_source_offset_buf;
  reg [33-1:0] _mul_37_rshift_source_size_buf;
  reg [32-1:0] _mul_37_rshift_source_stride_buf;
  reg [8-1:0] _mul_37_rshift_source_sel;
  reg [32-1:0] _mul_37_rshift_source_ram_raddr;
  reg _mul_37_rshift_source_ram_renable;
  wire [32-1:0] _mul_37_rshift_source_ram_rdata;
  reg _mul_37_rshift_source_fifo_deq;
  wire [32-1:0] _mul_37_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_37_rshift_source_empty_data;
  reg [33-1:0] _mul_37_z_sink_count;
  reg [5-1:0] _mul_37_z_sink_mode;
  reg [16-1:0] _mul_37_z_sink_generator_id;
  reg [32-1:0] _mul_37_z_sink_offset;
  reg [33-1:0] _mul_37_z_sink_size;
  reg [32-1:0] _mul_37_z_sink_stride;
  reg [32-1:0] _mul_37_z_sink_offset_buf;
  reg [33-1:0] _mul_37_z_sink_size_buf;
  reg [32-1:0] _mul_37_z_sink_stride_buf;
  reg [8-1:0] _mul_37_z_sink_sel;
  reg [32-1:0] _mul_37_z_sink_waddr;
  reg _mul_37_z_sink_wenable;
  reg [32-1:0] _mul_37_z_sink_wdata;
  reg _mul_37_z_sink_fifo_enq;
  reg [32-1:0] _mul_37_z_sink_fifo_wdata;
  reg [32-1:0] _mul_37_z_sink_immediate;
  reg _mul_38_stream_ivalid;
  wire _mul_38_stream_oready;
  wire _mul_38_stream_internal_oready;
  assign _mul_38_stream_internal_oready = 1;
  reg [32-1:0] _mul_38_fsm;
  localparam _mul_38_fsm_init = 0;
  wire _mul_38_run_flag;
  assign _mul_38_run_flag = 0;
  reg _mul_38_source_start;
  wire _mul_38_source_stop;
  reg _mul_38_source_busy;
  wire _mul_38_sink_start;
  wire _mul_38_sink_stop;
  wire _mul_38_sink_busy;
  wire _mul_38_busy;
  reg _mul_38_busy_reg;
  wire _mul_38_is_root;
  reg _mul_38_x_idle;
  reg [33-1:0] _mul_38_x_source_count;
  reg [5-1:0] _mul_38_x_source_mode;
  reg [16-1:0] _mul_38_x_source_generator_id;
  reg [32-1:0] _mul_38_x_source_offset;
  reg [33-1:0] _mul_38_x_source_size;
  reg [32-1:0] _mul_38_x_source_stride;
  reg [32-1:0] _mul_38_x_source_offset_buf;
  reg [33-1:0] _mul_38_x_source_size_buf;
  reg [32-1:0] _mul_38_x_source_stride_buf;
  reg [8-1:0] _mul_38_x_source_sel;
  reg [32-1:0] _mul_38_x_source_ram_raddr;
  reg _mul_38_x_source_ram_renable;
  wire [16-1:0] _mul_38_x_source_ram_rdata;
  reg _mul_38_x_source_fifo_deq;
  wire [16-1:0] _mul_38_x_source_fifo_rdata;
  reg [16-1:0] _mul_38_x_source_empty_data;
  reg _mul_38_y_idle;
  reg [33-1:0] _mul_38_y_source_count;
  reg [5-1:0] _mul_38_y_source_mode;
  reg [16-1:0] _mul_38_y_source_generator_id;
  reg [32-1:0] _mul_38_y_source_offset;
  reg [33-1:0] _mul_38_y_source_size;
  reg [32-1:0] _mul_38_y_source_stride;
  reg [32-1:0] _mul_38_y_source_offset_buf;
  reg [33-1:0] _mul_38_y_source_size_buf;
  reg [32-1:0] _mul_38_y_source_stride_buf;
  reg [8-1:0] _mul_38_y_source_sel;
  reg [32-1:0] _mul_38_y_source_ram_raddr;
  reg _mul_38_y_source_ram_renable;
  wire [16-1:0] _mul_38_y_source_ram_rdata;
  reg _mul_38_y_source_fifo_deq;
  wire [16-1:0] _mul_38_y_source_fifo_rdata;
  reg [16-1:0] _mul_38_y_source_empty_data;
  reg _mul_38_rshift_idle;
  reg [33-1:0] _mul_38_rshift_source_count;
  reg [5-1:0] _mul_38_rshift_source_mode;
  reg [16-1:0] _mul_38_rshift_source_generator_id;
  reg [32-1:0] _mul_38_rshift_source_offset;
  reg [33-1:0] _mul_38_rshift_source_size;
  reg [32-1:0] _mul_38_rshift_source_stride;
  reg [32-1:0] _mul_38_rshift_source_offset_buf;
  reg [33-1:0] _mul_38_rshift_source_size_buf;
  reg [32-1:0] _mul_38_rshift_source_stride_buf;
  reg [8-1:0] _mul_38_rshift_source_sel;
  reg [32-1:0] _mul_38_rshift_source_ram_raddr;
  reg _mul_38_rshift_source_ram_renable;
  wire [32-1:0] _mul_38_rshift_source_ram_rdata;
  reg _mul_38_rshift_source_fifo_deq;
  wire [32-1:0] _mul_38_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_38_rshift_source_empty_data;
  reg [33-1:0] _mul_38_z_sink_count;
  reg [5-1:0] _mul_38_z_sink_mode;
  reg [16-1:0] _mul_38_z_sink_generator_id;
  reg [32-1:0] _mul_38_z_sink_offset;
  reg [33-1:0] _mul_38_z_sink_size;
  reg [32-1:0] _mul_38_z_sink_stride;
  reg [32-1:0] _mul_38_z_sink_offset_buf;
  reg [33-1:0] _mul_38_z_sink_size_buf;
  reg [32-1:0] _mul_38_z_sink_stride_buf;
  reg [8-1:0] _mul_38_z_sink_sel;
  reg [32-1:0] _mul_38_z_sink_waddr;
  reg _mul_38_z_sink_wenable;
  reg [32-1:0] _mul_38_z_sink_wdata;
  reg _mul_38_z_sink_fifo_enq;
  reg [32-1:0] _mul_38_z_sink_fifo_wdata;
  reg [32-1:0] _mul_38_z_sink_immediate;
  reg _mul_39_stream_ivalid;
  wire _mul_39_stream_oready;
  wire _mul_39_stream_internal_oready;
  assign _mul_39_stream_internal_oready = 1;
  reg [32-1:0] _mul_39_fsm;
  localparam _mul_39_fsm_init = 0;
  wire _mul_39_run_flag;
  assign _mul_39_run_flag = 0;
  reg _mul_39_source_start;
  wire _mul_39_source_stop;
  reg _mul_39_source_busy;
  wire _mul_39_sink_start;
  wire _mul_39_sink_stop;
  wire _mul_39_sink_busy;
  wire _mul_39_busy;
  reg _mul_39_busy_reg;
  wire _mul_39_is_root;
  reg _mul_39_x_idle;
  reg [33-1:0] _mul_39_x_source_count;
  reg [5-1:0] _mul_39_x_source_mode;
  reg [16-1:0] _mul_39_x_source_generator_id;
  reg [32-1:0] _mul_39_x_source_offset;
  reg [33-1:0] _mul_39_x_source_size;
  reg [32-1:0] _mul_39_x_source_stride;
  reg [32-1:0] _mul_39_x_source_offset_buf;
  reg [33-1:0] _mul_39_x_source_size_buf;
  reg [32-1:0] _mul_39_x_source_stride_buf;
  reg [8-1:0] _mul_39_x_source_sel;
  reg [32-1:0] _mul_39_x_source_ram_raddr;
  reg _mul_39_x_source_ram_renable;
  wire [16-1:0] _mul_39_x_source_ram_rdata;
  reg _mul_39_x_source_fifo_deq;
  wire [16-1:0] _mul_39_x_source_fifo_rdata;
  reg [16-1:0] _mul_39_x_source_empty_data;
  reg _mul_39_y_idle;
  reg [33-1:0] _mul_39_y_source_count;
  reg [5-1:0] _mul_39_y_source_mode;
  reg [16-1:0] _mul_39_y_source_generator_id;
  reg [32-1:0] _mul_39_y_source_offset;
  reg [33-1:0] _mul_39_y_source_size;
  reg [32-1:0] _mul_39_y_source_stride;
  reg [32-1:0] _mul_39_y_source_offset_buf;
  reg [33-1:0] _mul_39_y_source_size_buf;
  reg [32-1:0] _mul_39_y_source_stride_buf;
  reg [8-1:0] _mul_39_y_source_sel;
  reg [32-1:0] _mul_39_y_source_ram_raddr;
  reg _mul_39_y_source_ram_renable;
  wire [16-1:0] _mul_39_y_source_ram_rdata;
  reg _mul_39_y_source_fifo_deq;
  wire [16-1:0] _mul_39_y_source_fifo_rdata;
  reg [16-1:0] _mul_39_y_source_empty_data;
  reg _mul_39_rshift_idle;
  reg [33-1:0] _mul_39_rshift_source_count;
  reg [5-1:0] _mul_39_rshift_source_mode;
  reg [16-1:0] _mul_39_rshift_source_generator_id;
  reg [32-1:0] _mul_39_rshift_source_offset;
  reg [33-1:0] _mul_39_rshift_source_size;
  reg [32-1:0] _mul_39_rshift_source_stride;
  reg [32-1:0] _mul_39_rshift_source_offset_buf;
  reg [33-1:0] _mul_39_rshift_source_size_buf;
  reg [32-1:0] _mul_39_rshift_source_stride_buf;
  reg [8-1:0] _mul_39_rshift_source_sel;
  reg [32-1:0] _mul_39_rshift_source_ram_raddr;
  reg _mul_39_rshift_source_ram_renable;
  wire [32-1:0] _mul_39_rshift_source_ram_rdata;
  reg _mul_39_rshift_source_fifo_deq;
  wire [32-1:0] _mul_39_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_39_rshift_source_empty_data;
  reg [33-1:0] _mul_39_z_sink_count;
  reg [5-1:0] _mul_39_z_sink_mode;
  reg [16-1:0] _mul_39_z_sink_generator_id;
  reg [32-1:0] _mul_39_z_sink_offset;
  reg [33-1:0] _mul_39_z_sink_size;
  reg [32-1:0] _mul_39_z_sink_stride;
  reg [32-1:0] _mul_39_z_sink_offset_buf;
  reg [33-1:0] _mul_39_z_sink_size_buf;
  reg [32-1:0] _mul_39_z_sink_stride_buf;
  reg [8-1:0] _mul_39_z_sink_sel;
  reg [32-1:0] _mul_39_z_sink_waddr;
  reg _mul_39_z_sink_wenable;
  reg [32-1:0] _mul_39_z_sink_wdata;
  reg _mul_39_z_sink_fifo_enq;
  reg [32-1:0] _mul_39_z_sink_fifo_wdata;
  reg [32-1:0] _mul_39_z_sink_immediate;
  reg _mul_40_stream_ivalid;
  wire _mul_40_stream_oready;
  wire _mul_40_stream_internal_oready;
  assign _mul_40_stream_internal_oready = 1;
  reg [32-1:0] _mul_40_fsm;
  localparam _mul_40_fsm_init = 0;
  wire _mul_40_run_flag;
  assign _mul_40_run_flag = 0;
  reg _mul_40_source_start;
  wire _mul_40_source_stop;
  reg _mul_40_source_busy;
  wire _mul_40_sink_start;
  wire _mul_40_sink_stop;
  wire _mul_40_sink_busy;
  wire _mul_40_busy;
  reg _mul_40_busy_reg;
  wire _mul_40_is_root;
  reg _mul_40_x_idle;
  reg [33-1:0] _mul_40_x_source_count;
  reg [5-1:0] _mul_40_x_source_mode;
  reg [16-1:0] _mul_40_x_source_generator_id;
  reg [32-1:0] _mul_40_x_source_offset;
  reg [33-1:0] _mul_40_x_source_size;
  reg [32-1:0] _mul_40_x_source_stride;
  reg [32-1:0] _mul_40_x_source_offset_buf;
  reg [33-1:0] _mul_40_x_source_size_buf;
  reg [32-1:0] _mul_40_x_source_stride_buf;
  reg [8-1:0] _mul_40_x_source_sel;
  reg [32-1:0] _mul_40_x_source_ram_raddr;
  reg _mul_40_x_source_ram_renable;
  wire [16-1:0] _mul_40_x_source_ram_rdata;
  reg _mul_40_x_source_fifo_deq;
  wire [16-1:0] _mul_40_x_source_fifo_rdata;
  reg [16-1:0] _mul_40_x_source_empty_data;
  reg _mul_40_y_idle;
  reg [33-1:0] _mul_40_y_source_count;
  reg [5-1:0] _mul_40_y_source_mode;
  reg [16-1:0] _mul_40_y_source_generator_id;
  reg [32-1:0] _mul_40_y_source_offset;
  reg [33-1:0] _mul_40_y_source_size;
  reg [32-1:0] _mul_40_y_source_stride;
  reg [32-1:0] _mul_40_y_source_offset_buf;
  reg [33-1:0] _mul_40_y_source_size_buf;
  reg [32-1:0] _mul_40_y_source_stride_buf;
  reg [8-1:0] _mul_40_y_source_sel;
  reg [32-1:0] _mul_40_y_source_ram_raddr;
  reg _mul_40_y_source_ram_renable;
  wire [16-1:0] _mul_40_y_source_ram_rdata;
  reg _mul_40_y_source_fifo_deq;
  wire [16-1:0] _mul_40_y_source_fifo_rdata;
  reg [16-1:0] _mul_40_y_source_empty_data;
  reg _mul_40_rshift_idle;
  reg [33-1:0] _mul_40_rshift_source_count;
  reg [5-1:0] _mul_40_rshift_source_mode;
  reg [16-1:0] _mul_40_rshift_source_generator_id;
  reg [32-1:0] _mul_40_rshift_source_offset;
  reg [33-1:0] _mul_40_rshift_source_size;
  reg [32-1:0] _mul_40_rshift_source_stride;
  reg [32-1:0] _mul_40_rshift_source_offset_buf;
  reg [33-1:0] _mul_40_rshift_source_size_buf;
  reg [32-1:0] _mul_40_rshift_source_stride_buf;
  reg [8-1:0] _mul_40_rshift_source_sel;
  reg [32-1:0] _mul_40_rshift_source_ram_raddr;
  reg _mul_40_rshift_source_ram_renable;
  wire [32-1:0] _mul_40_rshift_source_ram_rdata;
  reg _mul_40_rshift_source_fifo_deq;
  wire [32-1:0] _mul_40_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_40_rshift_source_empty_data;
  reg [33-1:0] _mul_40_z_sink_count;
  reg [5-1:0] _mul_40_z_sink_mode;
  reg [16-1:0] _mul_40_z_sink_generator_id;
  reg [32-1:0] _mul_40_z_sink_offset;
  reg [33-1:0] _mul_40_z_sink_size;
  reg [32-1:0] _mul_40_z_sink_stride;
  reg [32-1:0] _mul_40_z_sink_offset_buf;
  reg [33-1:0] _mul_40_z_sink_size_buf;
  reg [32-1:0] _mul_40_z_sink_stride_buf;
  reg [8-1:0] _mul_40_z_sink_sel;
  reg [32-1:0] _mul_40_z_sink_waddr;
  reg _mul_40_z_sink_wenable;
  reg [32-1:0] _mul_40_z_sink_wdata;
  reg _mul_40_z_sink_fifo_enq;
  reg [32-1:0] _mul_40_z_sink_fifo_wdata;
  reg [32-1:0] _mul_40_z_sink_immediate;
  reg _mul_41_stream_ivalid;
  wire _mul_41_stream_oready;
  wire _mul_41_stream_internal_oready;
  assign _mul_41_stream_internal_oready = 1;
  reg [32-1:0] _mul_41_fsm;
  localparam _mul_41_fsm_init = 0;
  wire _mul_41_run_flag;
  assign _mul_41_run_flag = 0;
  reg _mul_41_source_start;
  wire _mul_41_source_stop;
  reg _mul_41_source_busy;
  wire _mul_41_sink_start;
  wire _mul_41_sink_stop;
  wire _mul_41_sink_busy;
  wire _mul_41_busy;
  reg _mul_41_busy_reg;
  wire _mul_41_is_root;
  reg _mul_41_x_idle;
  reg [33-1:0] _mul_41_x_source_count;
  reg [5-1:0] _mul_41_x_source_mode;
  reg [16-1:0] _mul_41_x_source_generator_id;
  reg [32-1:0] _mul_41_x_source_offset;
  reg [33-1:0] _mul_41_x_source_size;
  reg [32-1:0] _mul_41_x_source_stride;
  reg [32-1:0] _mul_41_x_source_offset_buf;
  reg [33-1:0] _mul_41_x_source_size_buf;
  reg [32-1:0] _mul_41_x_source_stride_buf;
  reg [8-1:0] _mul_41_x_source_sel;
  reg [32-1:0] _mul_41_x_source_ram_raddr;
  reg _mul_41_x_source_ram_renable;
  wire [16-1:0] _mul_41_x_source_ram_rdata;
  reg _mul_41_x_source_fifo_deq;
  wire [16-1:0] _mul_41_x_source_fifo_rdata;
  reg [16-1:0] _mul_41_x_source_empty_data;
  reg _mul_41_y_idle;
  reg [33-1:0] _mul_41_y_source_count;
  reg [5-1:0] _mul_41_y_source_mode;
  reg [16-1:0] _mul_41_y_source_generator_id;
  reg [32-1:0] _mul_41_y_source_offset;
  reg [33-1:0] _mul_41_y_source_size;
  reg [32-1:0] _mul_41_y_source_stride;
  reg [32-1:0] _mul_41_y_source_offset_buf;
  reg [33-1:0] _mul_41_y_source_size_buf;
  reg [32-1:0] _mul_41_y_source_stride_buf;
  reg [8-1:0] _mul_41_y_source_sel;
  reg [32-1:0] _mul_41_y_source_ram_raddr;
  reg _mul_41_y_source_ram_renable;
  wire [16-1:0] _mul_41_y_source_ram_rdata;
  reg _mul_41_y_source_fifo_deq;
  wire [16-1:0] _mul_41_y_source_fifo_rdata;
  reg [16-1:0] _mul_41_y_source_empty_data;
  reg _mul_41_rshift_idle;
  reg [33-1:0] _mul_41_rshift_source_count;
  reg [5-1:0] _mul_41_rshift_source_mode;
  reg [16-1:0] _mul_41_rshift_source_generator_id;
  reg [32-1:0] _mul_41_rshift_source_offset;
  reg [33-1:0] _mul_41_rshift_source_size;
  reg [32-1:0] _mul_41_rshift_source_stride;
  reg [32-1:0] _mul_41_rshift_source_offset_buf;
  reg [33-1:0] _mul_41_rshift_source_size_buf;
  reg [32-1:0] _mul_41_rshift_source_stride_buf;
  reg [8-1:0] _mul_41_rshift_source_sel;
  reg [32-1:0] _mul_41_rshift_source_ram_raddr;
  reg _mul_41_rshift_source_ram_renable;
  wire [32-1:0] _mul_41_rshift_source_ram_rdata;
  reg _mul_41_rshift_source_fifo_deq;
  wire [32-1:0] _mul_41_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_41_rshift_source_empty_data;
  reg [33-1:0] _mul_41_z_sink_count;
  reg [5-1:0] _mul_41_z_sink_mode;
  reg [16-1:0] _mul_41_z_sink_generator_id;
  reg [32-1:0] _mul_41_z_sink_offset;
  reg [33-1:0] _mul_41_z_sink_size;
  reg [32-1:0] _mul_41_z_sink_stride;
  reg [32-1:0] _mul_41_z_sink_offset_buf;
  reg [33-1:0] _mul_41_z_sink_size_buf;
  reg [32-1:0] _mul_41_z_sink_stride_buf;
  reg [8-1:0] _mul_41_z_sink_sel;
  reg [32-1:0] _mul_41_z_sink_waddr;
  reg _mul_41_z_sink_wenable;
  reg [32-1:0] _mul_41_z_sink_wdata;
  reg _mul_41_z_sink_fifo_enq;
  reg [32-1:0] _mul_41_z_sink_fifo_wdata;
  reg [32-1:0] _mul_41_z_sink_immediate;
  reg _mul_42_stream_ivalid;
  wire _mul_42_stream_oready;
  wire _mul_42_stream_internal_oready;
  assign _mul_42_stream_internal_oready = 1;
  reg [32-1:0] _mul_42_fsm;
  localparam _mul_42_fsm_init = 0;
  wire _mul_42_run_flag;
  assign _mul_42_run_flag = 0;
  reg _mul_42_source_start;
  wire _mul_42_source_stop;
  reg _mul_42_source_busy;
  wire _mul_42_sink_start;
  wire _mul_42_sink_stop;
  wire _mul_42_sink_busy;
  wire _mul_42_busy;
  reg _mul_42_busy_reg;
  wire _mul_42_is_root;
  reg _mul_42_x_idle;
  reg [33-1:0] _mul_42_x_source_count;
  reg [5-1:0] _mul_42_x_source_mode;
  reg [16-1:0] _mul_42_x_source_generator_id;
  reg [32-1:0] _mul_42_x_source_offset;
  reg [33-1:0] _mul_42_x_source_size;
  reg [32-1:0] _mul_42_x_source_stride;
  reg [32-1:0] _mul_42_x_source_offset_buf;
  reg [33-1:0] _mul_42_x_source_size_buf;
  reg [32-1:0] _mul_42_x_source_stride_buf;
  reg [8-1:0] _mul_42_x_source_sel;
  reg [32-1:0] _mul_42_x_source_ram_raddr;
  reg _mul_42_x_source_ram_renable;
  wire [16-1:0] _mul_42_x_source_ram_rdata;
  reg _mul_42_x_source_fifo_deq;
  wire [16-1:0] _mul_42_x_source_fifo_rdata;
  reg [16-1:0] _mul_42_x_source_empty_data;
  reg _mul_42_y_idle;
  reg [33-1:0] _mul_42_y_source_count;
  reg [5-1:0] _mul_42_y_source_mode;
  reg [16-1:0] _mul_42_y_source_generator_id;
  reg [32-1:0] _mul_42_y_source_offset;
  reg [33-1:0] _mul_42_y_source_size;
  reg [32-1:0] _mul_42_y_source_stride;
  reg [32-1:0] _mul_42_y_source_offset_buf;
  reg [33-1:0] _mul_42_y_source_size_buf;
  reg [32-1:0] _mul_42_y_source_stride_buf;
  reg [8-1:0] _mul_42_y_source_sel;
  reg [32-1:0] _mul_42_y_source_ram_raddr;
  reg _mul_42_y_source_ram_renable;
  wire [16-1:0] _mul_42_y_source_ram_rdata;
  reg _mul_42_y_source_fifo_deq;
  wire [16-1:0] _mul_42_y_source_fifo_rdata;
  reg [16-1:0] _mul_42_y_source_empty_data;
  reg _mul_42_rshift_idle;
  reg [33-1:0] _mul_42_rshift_source_count;
  reg [5-1:0] _mul_42_rshift_source_mode;
  reg [16-1:0] _mul_42_rshift_source_generator_id;
  reg [32-1:0] _mul_42_rshift_source_offset;
  reg [33-1:0] _mul_42_rshift_source_size;
  reg [32-1:0] _mul_42_rshift_source_stride;
  reg [32-1:0] _mul_42_rshift_source_offset_buf;
  reg [33-1:0] _mul_42_rshift_source_size_buf;
  reg [32-1:0] _mul_42_rshift_source_stride_buf;
  reg [8-1:0] _mul_42_rshift_source_sel;
  reg [32-1:0] _mul_42_rshift_source_ram_raddr;
  reg _mul_42_rshift_source_ram_renable;
  wire [32-1:0] _mul_42_rshift_source_ram_rdata;
  reg _mul_42_rshift_source_fifo_deq;
  wire [32-1:0] _mul_42_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_42_rshift_source_empty_data;
  reg [33-1:0] _mul_42_z_sink_count;
  reg [5-1:0] _mul_42_z_sink_mode;
  reg [16-1:0] _mul_42_z_sink_generator_id;
  reg [32-1:0] _mul_42_z_sink_offset;
  reg [33-1:0] _mul_42_z_sink_size;
  reg [32-1:0] _mul_42_z_sink_stride;
  reg [32-1:0] _mul_42_z_sink_offset_buf;
  reg [33-1:0] _mul_42_z_sink_size_buf;
  reg [32-1:0] _mul_42_z_sink_stride_buf;
  reg [8-1:0] _mul_42_z_sink_sel;
  reg [32-1:0] _mul_42_z_sink_waddr;
  reg _mul_42_z_sink_wenable;
  reg [32-1:0] _mul_42_z_sink_wdata;
  reg _mul_42_z_sink_fifo_enq;
  reg [32-1:0] _mul_42_z_sink_fifo_wdata;
  reg [32-1:0] _mul_42_z_sink_immediate;
  reg _mul_43_stream_ivalid;
  wire _mul_43_stream_oready;
  wire _mul_43_stream_internal_oready;
  assign _mul_43_stream_internal_oready = 1;
  reg [32-1:0] _mul_43_fsm;
  localparam _mul_43_fsm_init = 0;
  wire _mul_43_run_flag;
  assign _mul_43_run_flag = 0;
  reg _mul_43_source_start;
  wire _mul_43_source_stop;
  reg _mul_43_source_busy;
  wire _mul_43_sink_start;
  wire _mul_43_sink_stop;
  wire _mul_43_sink_busy;
  wire _mul_43_busy;
  reg _mul_43_busy_reg;
  wire _mul_43_is_root;
  reg _mul_43_x_idle;
  reg [33-1:0] _mul_43_x_source_count;
  reg [5-1:0] _mul_43_x_source_mode;
  reg [16-1:0] _mul_43_x_source_generator_id;
  reg [32-1:0] _mul_43_x_source_offset;
  reg [33-1:0] _mul_43_x_source_size;
  reg [32-1:0] _mul_43_x_source_stride;
  reg [32-1:0] _mul_43_x_source_offset_buf;
  reg [33-1:0] _mul_43_x_source_size_buf;
  reg [32-1:0] _mul_43_x_source_stride_buf;
  reg [8-1:0] _mul_43_x_source_sel;
  reg [32-1:0] _mul_43_x_source_ram_raddr;
  reg _mul_43_x_source_ram_renable;
  wire [16-1:0] _mul_43_x_source_ram_rdata;
  reg _mul_43_x_source_fifo_deq;
  wire [16-1:0] _mul_43_x_source_fifo_rdata;
  reg [16-1:0] _mul_43_x_source_empty_data;
  reg _mul_43_y_idle;
  reg [33-1:0] _mul_43_y_source_count;
  reg [5-1:0] _mul_43_y_source_mode;
  reg [16-1:0] _mul_43_y_source_generator_id;
  reg [32-1:0] _mul_43_y_source_offset;
  reg [33-1:0] _mul_43_y_source_size;
  reg [32-1:0] _mul_43_y_source_stride;
  reg [32-1:0] _mul_43_y_source_offset_buf;
  reg [33-1:0] _mul_43_y_source_size_buf;
  reg [32-1:0] _mul_43_y_source_stride_buf;
  reg [8-1:0] _mul_43_y_source_sel;
  reg [32-1:0] _mul_43_y_source_ram_raddr;
  reg _mul_43_y_source_ram_renable;
  wire [16-1:0] _mul_43_y_source_ram_rdata;
  reg _mul_43_y_source_fifo_deq;
  wire [16-1:0] _mul_43_y_source_fifo_rdata;
  reg [16-1:0] _mul_43_y_source_empty_data;
  reg _mul_43_rshift_idle;
  reg [33-1:0] _mul_43_rshift_source_count;
  reg [5-1:0] _mul_43_rshift_source_mode;
  reg [16-1:0] _mul_43_rshift_source_generator_id;
  reg [32-1:0] _mul_43_rshift_source_offset;
  reg [33-1:0] _mul_43_rshift_source_size;
  reg [32-1:0] _mul_43_rshift_source_stride;
  reg [32-1:0] _mul_43_rshift_source_offset_buf;
  reg [33-1:0] _mul_43_rshift_source_size_buf;
  reg [32-1:0] _mul_43_rshift_source_stride_buf;
  reg [8-1:0] _mul_43_rshift_source_sel;
  reg [32-1:0] _mul_43_rshift_source_ram_raddr;
  reg _mul_43_rshift_source_ram_renable;
  wire [32-1:0] _mul_43_rshift_source_ram_rdata;
  reg _mul_43_rshift_source_fifo_deq;
  wire [32-1:0] _mul_43_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_43_rshift_source_empty_data;
  reg [33-1:0] _mul_43_z_sink_count;
  reg [5-1:0] _mul_43_z_sink_mode;
  reg [16-1:0] _mul_43_z_sink_generator_id;
  reg [32-1:0] _mul_43_z_sink_offset;
  reg [33-1:0] _mul_43_z_sink_size;
  reg [32-1:0] _mul_43_z_sink_stride;
  reg [32-1:0] _mul_43_z_sink_offset_buf;
  reg [33-1:0] _mul_43_z_sink_size_buf;
  reg [32-1:0] _mul_43_z_sink_stride_buf;
  reg [8-1:0] _mul_43_z_sink_sel;
  reg [32-1:0] _mul_43_z_sink_waddr;
  reg _mul_43_z_sink_wenable;
  reg [32-1:0] _mul_43_z_sink_wdata;
  reg _mul_43_z_sink_fifo_enq;
  reg [32-1:0] _mul_43_z_sink_fifo_wdata;
  reg [32-1:0] _mul_43_z_sink_immediate;
  reg __reduce_max_44_stream_ivalid;
  wire __reduce_max_44_stream_oready;
  wire __reduce_max_44_stream_internal_oready;
  assign __reduce_max_44_stream_internal_oready = 1;
  reg [32-1:0] __reduce_max_44_fsm;
  localparam __reduce_max_44_fsm_init = 0;
  wire __reduce_max_44_run_flag;
  assign __reduce_max_44_run_flag = 0;
  reg __reduce_max_44_source_start;
  wire __reduce_max_44_source_stop;
  reg __reduce_max_44_source_busy;
  wire __reduce_max_44_sink_start;
  wire __reduce_max_44_sink_stop;
  wire __reduce_max_44_sink_busy;
  wire __reduce_max_44_busy;
  reg __reduce_max_44_busy_reg;
  wire __reduce_max_44_is_root;
  reg __reduce_max_44_x_idle;
  reg [33-1:0] __reduce_max_44_x_source_count;
  reg [5-1:0] __reduce_max_44_x_source_mode;
  reg [16-1:0] __reduce_max_44_x_source_generator_id;
  reg [32-1:0] __reduce_max_44_x_source_offset;
  reg [33-1:0] __reduce_max_44_x_source_size;
  reg [32-1:0] __reduce_max_44_x_source_stride;
  reg [32-1:0] __reduce_max_44_x_source_offset_buf;
  reg [33-1:0] __reduce_max_44_x_source_size_buf;
  reg [32-1:0] __reduce_max_44_x_source_stride_buf;
  reg [8-1:0] __reduce_max_44_x_source_sel;
  reg [32-1:0] __reduce_max_44_x_source_ram_raddr;
  reg __reduce_max_44_x_source_ram_renable;
  wire [16-1:0] __reduce_max_44_x_source_ram_rdata;
  reg __reduce_max_44_x_source_fifo_deq;
  wire [16-1:0] __reduce_max_44_x_source_fifo_rdata;
  reg [16-1:0] __reduce_max_44_x_source_empty_data;
  reg [32-1:0] __reduce_max_44_size_next_parameter_data;
  reg [33-1:0] __reduce_max_44_data_sink_count;
  reg [5-1:0] __reduce_max_44_data_sink_mode;
  reg [16-1:0] __reduce_max_44_data_sink_generator_id;
  reg [32-1:0] __reduce_max_44_data_sink_offset;
  reg [33-1:0] __reduce_max_44_data_sink_size;
  reg [32-1:0] __reduce_max_44_data_sink_stride;
  reg [32-1:0] __reduce_max_44_data_sink_offset_buf;
  reg [33-1:0] __reduce_max_44_data_sink_size_buf;
  reg [32-1:0] __reduce_max_44_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_44_data_sink_sel;
  reg [32-1:0] __reduce_max_44_data_sink_waddr;
  reg __reduce_max_44_data_sink_wenable;
  reg [16-1:0] __reduce_max_44_data_sink_wdata;
  reg __reduce_max_44_data_sink_fifo_enq;
  reg [16-1:0] __reduce_max_44_data_sink_fifo_wdata;
  reg [16-1:0] __reduce_max_44_data_sink_immediate;
  reg [33-1:0] __reduce_max_44_valid_sink_count;
  reg [5-1:0] __reduce_max_44_valid_sink_mode;
  reg [16-1:0] __reduce_max_44_valid_sink_generator_id;
  reg [32-1:0] __reduce_max_44_valid_sink_offset;
  reg [33-1:0] __reduce_max_44_valid_sink_size;
  reg [32-1:0] __reduce_max_44_valid_sink_stride;
  reg [32-1:0] __reduce_max_44_valid_sink_offset_buf;
  reg [33-1:0] __reduce_max_44_valid_sink_size_buf;
  reg [32-1:0] __reduce_max_44_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_44_valid_sink_sel;
  reg [32-1:0] __reduce_max_44_valid_sink_waddr;
  reg __reduce_max_44_valid_sink_wenable;
  reg [1-1:0] __reduce_max_44_valid_sink_wdata;
  reg __reduce_max_44_valid_sink_fifo_enq;
  reg [1-1:0] __reduce_max_44_valid_sink_fifo_wdata;
  reg [1-1:0] __reduce_max_44_valid_sink_immediate;
  reg __reduce_max_45_stream_ivalid;
  wire __reduce_max_45_stream_oready;
  wire __reduce_max_45_stream_internal_oready;
  assign __reduce_max_45_stream_internal_oready = 1;
  reg [32-1:0] __reduce_max_45_fsm;
  localparam __reduce_max_45_fsm_init = 0;
  wire __reduce_max_45_run_flag;
  assign __reduce_max_45_run_flag = 0;
  reg __reduce_max_45_source_start;
  wire __reduce_max_45_source_stop;
  reg __reduce_max_45_source_busy;
  wire __reduce_max_45_sink_start;
  wire __reduce_max_45_sink_stop;
  wire __reduce_max_45_sink_busy;
  wire __reduce_max_45_busy;
  reg __reduce_max_45_busy_reg;
  wire __reduce_max_45_is_root;
  reg __reduce_max_45_x_idle;
  reg [33-1:0] __reduce_max_45_x_source_count;
  reg [5-1:0] __reduce_max_45_x_source_mode;
  reg [16-1:0] __reduce_max_45_x_source_generator_id;
  reg [32-1:0] __reduce_max_45_x_source_offset;
  reg [33-1:0] __reduce_max_45_x_source_size;
  reg [32-1:0] __reduce_max_45_x_source_stride;
  reg [32-1:0] __reduce_max_45_x_source_offset_buf;
  reg [33-1:0] __reduce_max_45_x_source_size_buf;
  reg [32-1:0] __reduce_max_45_x_source_stride_buf;
  reg [8-1:0] __reduce_max_45_x_source_sel;
  reg [32-1:0] __reduce_max_45_x_source_ram_raddr;
  reg __reduce_max_45_x_source_ram_renable;
  wire [16-1:0] __reduce_max_45_x_source_ram_rdata;
  reg __reduce_max_45_x_source_fifo_deq;
  wire [16-1:0] __reduce_max_45_x_source_fifo_rdata;
  reg [16-1:0] __reduce_max_45_x_source_empty_data;
  reg [32-1:0] __reduce_max_45_size_next_parameter_data;
  reg [33-1:0] __reduce_max_45_data_sink_count;
  reg [5-1:0] __reduce_max_45_data_sink_mode;
  reg [16-1:0] __reduce_max_45_data_sink_generator_id;
  reg [32-1:0] __reduce_max_45_data_sink_offset;
  reg [33-1:0] __reduce_max_45_data_sink_size;
  reg [32-1:0] __reduce_max_45_data_sink_stride;
  reg [32-1:0] __reduce_max_45_data_sink_offset_buf;
  reg [33-1:0] __reduce_max_45_data_sink_size_buf;
  reg [32-1:0] __reduce_max_45_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_45_data_sink_sel;
  reg [32-1:0] __reduce_max_45_data_sink_waddr;
  reg __reduce_max_45_data_sink_wenable;
  reg [16-1:0] __reduce_max_45_data_sink_wdata;
  reg __reduce_max_45_data_sink_fifo_enq;
  reg [16-1:0] __reduce_max_45_data_sink_fifo_wdata;
  reg [16-1:0] __reduce_max_45_data_sink_immediate;
  reg [33-1:0] __reduce_max_45_valid_sink_count;
  reg [5-1:0] __reduce_max_45_valid_sink_mode;
  reg [16-1:0] __reduce_max_45_valid_sink_generator_id;
  reg [32-1:0] __reduce_max_45_valid_sink_offset;
  reg [33-1:0] __reduce_max_45_valid_sink_size;
  reg [32-1:0] __reduce_max_45_valid_sink_stride;
  reg [32-1:0] __reduce_max_45_valid_sink_offset_buf;
  reg [33-1:0] __reduce_max_45_valid_sink_size_buf;
  reg [32-1:0] __reduce_max_45_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_45_valid_sink_sel;
  reg [32-1:0] __reduce_max_45_valid_sink_waddr;
  reg __reduce_max_45_valid_sink_wenable;
  reg [1-1:0] __reduce_max_45_valid_sink_wdata;
  reg __reduce_max_45_valid_sink_fifo_enq;
  reg [1-1:0] __reduce_max_45_valid_sink_fifo_wdata;
  reg [1-1:0] __reduce_max_45_valid_sink_immediate;
  reg _stream_conv2d_4_stream_ivalid;
  wire _stream_conv2d_4_stream_oready;
  wire _stream_conv2d_4_stream_internal_oready;
  assign _stream_conv2d_4_stream_oready = _stream_conv2d_4_stream_internal_oready;
  reg [32-1:0] _stream_conv2d_4_fsm;
  localparam _stream_conv2d_4_fsm_init = 0;
  wire _stream_conv2d_4_run_flag;
  reg _stream_conv2d_4_source_start;
  wire _stream_conv2d_4_source_stop;
  reg _stream_conv2d_4_source_busy;
  wire _stream_conv2d_4_sink_start;
  wire _stream_conv2d_4_sink_stop;
  wire _stream_conv2d_4_sink_busy;
  wire _stream_conv2d_4_busy;
  reg _stream_conv2d_4_busy_reg;
  wire _stream_conv2d_4_is_root;
  assign _stream_conv2d_4_is_root = 1;
  reg [6-1:0] _stream_conv2d_4_parameter_0_next_parameter_data;
  reg [2-1:0] _stream_conv2d_4_parameter_1_next_parameter_data;
  reg [2-1:0] _stream_conv2d_4_parameter_2_next_parameter_data;
  reg [9-1:0] _stream_conv2d_4_parameter_3_next_parameter_data;
  reg [2-1:0] _stream_conv2d_4_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_6_next_parameter_data;
  reg _stream_conv2d_4_source_7_idle;
  reg [33-1:0] _stream_conv2d_4_source_7_source_count;
  reg [5-1:0] _stream_conv2d_4_source_7_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_7_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_7_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_7_source_size;
  reg [32-1:0] _stream_conv2d_4_source_7_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_7_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_7_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_7_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_7_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_7_source_ram_raddr;
  reg _stream_conv2d_4_source_7_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_7_source_ram_rdata;
  reg _stream_conv2d_4_source_7_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_7_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_7_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_8_next_parameter_data;
  reg _stream_conv2d_4_source_9_idle;
  reg [33-1:0] _stream_conv2d_4_source_9_source_count;
  reg [5-1:0] _stream_conv2d_4_source_9_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_9_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_9_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_9_source_size;
  reg [32-1:0] _stream_conv2d_4_source_9_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_9_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_9_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_9_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_9_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_9_source_ram_raddr;
  reg _stream_conv2d_4_source_9_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_9_source_ram_rdata;
  reg _stream_conv2d_4_source_9_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_9_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_9_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_10_next_parameter_data;
  reg _stream_conv2d_4_source_11_idle;
  reg [33-1:0] _stream_conv2d_4_source_11_source_count;
  reg [5-1:0] _stream_conv2d_4_source_11_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_11_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_11_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_11_source_size;
  reg [32-1:0] _stream_conv2d_4_source_11_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_11_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_11_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_11_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_11_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_11_source_ram_raddr;
  reg _stream_conv2d_4_source_11_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_11_source_ram_rdata;
  reg _stream_conv2d_4_source_11_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_11_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_11_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_12_next_parameter_data;
  reg _stream_conv2d_4_source_13_idle;
  reg [33-1:0] _stream_conv2d_4_source_13_source_count;
  reg [5-1:0] _stream_conv2d_4_source_13_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_13_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_13_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_13_source_size;
  reg [32-1:0] _stream_conv2d_4_source_13_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_13_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_13_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_13_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_13_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_13_source_ram_raddr;
  reg _stream_conv2d_4_source_13_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_13_source_ram_rdata;
  reg _stream_conv2d_4_source_13_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_13_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_13_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_14_next_parameter_data;
  reg _stream_conv2d_4_source_15_idle;
  reg [33-1:0] _stream_conv2d_4_source_15_source_count;
  reg [5-1:0] _stream_conv2d_4_source_15_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_15_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_15_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_15_source_size;
  reg [32-1:0] _stream_conv2d_4_source_15_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_15_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_15_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_15_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_15_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_15_source_ram_raddr;
  reg _stream_conv2d_4_source_15_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_15_source_ram_rdata;
  reg _stream_conv2d_4_source_15_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_15_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_15_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_conv2d_4_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_19_next_parameter_data;
  reg _stream_conv2d_4_source_20_idle;
  reg [33-1:0] _stream_conv2d_4_source_20_source_count;
  reg [5-1:0] _stream_conv2d_4_source_20_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_20_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_20_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_20_source_size;
  reg [32-1:0] _stream_conv2d_4_source_20_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_20_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_20_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_20_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_20_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_20_source_ram_raddr;
  reg _stream_conv2d_4_source_20_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_20_source_ram_rdata;
  reg _stream_conv2d_4_source_20_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_20_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_20_source_empty_data;
  reg _stream_conv2d_4_source_21_idle;
  reg [33-1:0] _stream_conv2d_4_source_21_source_count;
  reg [5-1:0] _stream_conv2d_4_source_21_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_21_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_21_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_21_source_size;
  reg [32-1:0] _stream_conv2d_4_source_21_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_21_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_21_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_21_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_21_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_21_source_ram_raddr;
  reg _stream_conv2d_4_source_21_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_21_source_ram_rdata;
  reg _stream_conv2d_4_source_21_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_21_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_21_source_empty_data;
  reg _stream_conv2d_4_source_22_idle;
  reg [33-1:0] _stream_conv2d_4_source_22_source_count;
  reg [5-1:0] _stream_conv2d_4_source_22_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_22_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_22_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_22_source_size;
  reg [32-1:0] _stream_conv2d_4_source_22_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_22_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_22_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_22_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_22_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_22_source_ram_raddr;
  reg _stream_conv2d_4_source_22_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_22_source_ram_rdata;
  reg _stream_conv2d_4_source_22_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_22_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_22_source_empty_data;
  reg _stream_conv2d_4_source_23_idle;
  reg [33-1:0] _stream_conv2d_4_source_23_source_count;
  reg [5-1:0] _stream_conv2d_4_source_23_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_23_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_23_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_23_source_size;
  reg [32-1:0] _stream_conv2d_4_source_23_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_23_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_23_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_23_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_23_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_23_source_ram_raddr;
  reg _stream_conv2d_4_source_23_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_23_source_ram_rdata;
  reg _stream_conv2d_4_source_23_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_23_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_23_source_empty_data;
  reg _stream_conv2d_4_source_24_idle;
  reg [33-1:0] _stream_conv2d_4_source_24_source_count;
  reg [5-1:0] _stream_conv2d_4_source_24_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_24_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_24_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_24_source_size;
  reg [32-1:0] _stream_conv2d_4_source_24_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_24_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_24_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_24_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_24_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_24_source_ram_raddr;
  reg _stream_conv2d_4_source_24_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_24_source_ram_rdata;
  reg _stream_conv2d_4_source_24_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_24_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_24_source_empty_data;
  reg _stream_conv2d_4_source_25_idle;
  reg [33-1:0] _stream_conv2d_4_source_25_source_count;
  reg [5-1:0] _stream_conv2d_4_source_25_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_25_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_25_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_25_source_size;
  reg [32-1:0] _stream_conv2d_4_source_25_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_25_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_25_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_25_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_25_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_25_source_ram_raddr;
  reg _stream_conv2d_4_source_25_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_25_source_ram_rdata;
  reg _stream_conv2d_4_source_25_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_25_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_25_source_empty_data;
  reg _stream_conv2d_4_source_26_idle;
  reg [33-1:0] _stream_conv2d_4_source_26_source_count;
  reg [5-1:0] _stream_conv2d_4_source_26_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_26_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_26_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_26_source_size;
  reg [32-1:0] _stream_conv2d_4_source_26_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_26_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_26_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_26_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_26_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_26_source_ram_raddr;
  reg _stream_conv2d_4_source_26_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_26_source_ram_rdata;
  reg _stream_conv2d_4_source_26_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_26_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_26_source_empty_data;
  reg _stream_conv2d_4_source_27_idle;
  reg [33-1:0] _stream_conv2d_4_source_27_source_count;
  reg [5-1:0] _stream_conv2d_4_source_27_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_27_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_27_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_27_source_size;
  reg [32-1:0] _stream_conv2d_4_source_27_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_27_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_27_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_27_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_27_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_27_source_ram_raddr;
  reg _stream_conv2d_4_source_27_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_27_source_ram_rdata;
  reg _stream_conv2d_4_source_27_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_27_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_27_source_empty_data;
  reg _stream_conv2d_4_source_28_idle;
  reg [33-1:0] _stream_conv2d_4_source_28_source_count;
  reg [5-1:0] _stream_conv2d_4_source_28_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_28_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_28_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_28_source_size;
  reg [32-1:0] _stream_conv2d_4_source_28_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_28_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_28_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_28_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_28_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_28_source_ram_raddr;
  reg _stream_conv2d_4_source_28_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_28_source_ram_rdata;
  reg _stream_conv2d_4_source_28_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_28_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_28_source_empty_data;
  reg _stream_conv2d_4_source_29_idle;
  reg [33-1:0] _stream_conv2d_4_source_29_source_count;
  reg [5-1:0] _stream_conv2d_4_source_29_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_29_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_29_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_29_source_size;
  reg [32-1:0] _stream_conv2d_4_source_29_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_29_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_29_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_29_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_29_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_29_source_ram_raddr;
  reg _stream_conv2d_4_source_29_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_29_source_ram_rdata;
  reg _stream_conv2d_4_source_29_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_29_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_29_source_empty_data;
  reg _stream_conv2d_4_source_30_idle;
  reg [33-1:0] _stream_conv2d_4_source_30_source_count;
  reg [5-1:0] _stream_conv2d_4_source_30_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_30_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_30_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_30_source_size;
  reg [32-1:0] _stream_conv2d_4_source_30_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_30_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_30_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_30_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_30_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_30_source_ram_raddr;
  reg _stream_conv2d_4_source_30_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_30_source_ram_rdata;
  reg _stream_conv2d_4_source_30_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_30_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_30_source_empty_data;
  reg _stream_conv2d_4_source_31_idle;
  reg [33-1:0] _stream_conv2d_4_source_31_source_count;
  reg [5-1:0] _stream_conv2d_4_source_31_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_31_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_31_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_31_source_size;
  reg [32-1:0] _stream_conv2d_4_source_31_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_31_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_31_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_31_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_31_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_31_source_ram_raddr;
  reg _stream_conv2d_4_source_31_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_31_source_ram_rdata;
  reg _stream_conv2d_4_source_31_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_31_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_31_source_empty_data;
  reg _stream_conv2d_4_source_32_idle;
  reg [33-1:0] _stream_conv2d_4_source_32_source_count;
  reg [5-1:0] _stream_conv2d_4_source_32_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_32_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_32_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_32_source_size;
  reg [32-1:0] _stream_conv2d_4_source_32_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_32_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_32_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_32_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_32_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_32_source_ram_raddr;
  reg _stream_conv2d_4_source_32_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_32_source_ram_rdata;
  reg _stream_conv2d_4_source_32_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_32_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_32_source_empty_data;
  reg _stream_conv2d_4_source_33_idle;
  reg [33-1:0] _stream_conv2d_4_source_33_source_count;
  reg [5-1:0] _stream_conv2d_4_source_33_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_33_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_33_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_33_source_size;
  reg [32-1:0] _stream_conv2d_4_source_33_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_33_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_33_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_33_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_33_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_33_source_ram_raddr;
  reg _stream_conv2d_4_source_33_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_33_source_ram_rdata;
  reg _stream_conv2d_4_source_33_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_33_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_33_source_empty_data;
  reg _stream_conv2d_4_source_34_idle;
  reg [33-1:0] _stream_conv2d_4_source_34_source_count;
  reg [5-1:0] _stream_conv2d_4_source_34_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_34_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_34_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_34_source_size;
  reg [32-1:0] _stream_conv2d_4_source_34_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_34_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_34_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_34_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_34_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_34_source_ram_raddr;
  reg _stream_conv2d_4_source_34_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_34_source_ram_rdata;
  reg _stream_conv2d_4_source_34_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_34_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_34_source_empty_data;
  reg _stream_conv2d_4_source_35_idle;
  reg [33-1:0] _stream_conv2d_4_source_35_source_count;
  reg [5-1:0] _stream_conv2d_4_source_35_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_35_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_35_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_35_source_size;
  reg [32-1:0] _stream_conv2d_4_source_35_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_35_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_35_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_35_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_35_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_35_source_ram_raddr;
  reg _stream_conv2d_4_source_35_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_35_source_ram_rdata;
  reg _stream_conv2d_4_source_35_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_35_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_35_source_empty_data;
  reg _stream_conv2d_4_source_36_idle;
  reg [33-1:0] _stream_conv2d_4_source_36_source_count;
  reg [5-1:0] _stream_conv2d_4_source_36_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_36_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_36_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_36_source_size;
  reg [32-1:0] _stream_conv2d_4_source_36_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_36_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_36_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_36_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_36_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_36_source_ram_raddr;
  reg _stream_conv2d_4_source_36_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_36_source_ram_rdata;
  reg _stream_conv2d_4_source_36_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_36_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_36_source_empty_data;
  reg _stream_conv2d_4_source_37_idle;
  reg [33-1:0] _stream_conv2d_4_source_37_source_count;
  reg [5-1:0] _stream_conv2d_4_source_37_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_37_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_37_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_37_source_size;
  reg [32-1:0] _stream_conv2d_4_source_37_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_37_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_37_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_37_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_37_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_37_source_ram_raddr;
  reg _stream_conv2d_4_source_37_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_37_source_ram_rdata;
  reg _stream_conv2d_4_source_37_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_37_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_37_source_empty_data;
  reg _stream_conv2d_4_source_38_idle;
  reg [33-1:0] _stream_conv2d_4_source_38_source_count;
  reg [5-1:0] _stream_conv2d_4_source_38_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_38_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_38_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_38_source_size;
  reg [32-1:0] _stream_conv2d_4_source_38_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_38_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_38_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_38_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_38_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_38_source_ram_raddr;
  reg _stream_conv2d_4_source_38_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_38_source_ram_rdata;
  reg _stream_conv2d_4_source_38_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_38_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_38_source_empty_data;
  reg _stream_conv2d_4_source_39_idle;
  reg [33-1:0] _stream_conv2d_4_source_39_source_count;
  reg [5-1:0] _stream_conv2d_4_source_39_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_39_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_39_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_39_source_size;
  reg [32-1:0] _stream_conv2d_4_source_39_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_39_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_39_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_39_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_39_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_39_source_ram_raddr;
  reg _stream_conv2d_4_source_39_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_39_source_ram_rdata;
  reg _stream_conv2d_4_source_39_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_39_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_39_source_empty_data;
  reg _stream_conv2d_4_source_40_idle;
  reg [33-1:0] _stream_conv2d_4_source_40_source_count;
  reg [5-1:0] _stream_conv2d_4_source_40_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_40_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_40_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_40_source_size;
  reg [32-1:0] _stream_conv2d_4_source_40_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_40_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_40_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_40_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_40_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_40_source_ram_raddr;
  reg _stream_conv2d_4_source_40_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_40_source_ram_rdata;
  reg _stream_conv2d_4_source_40_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_40_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_40_source_empty_data;
  reg _stream_conv2d_4_source_41_idle;
  reg [33-1:0] _stream_conv2d_4_source_41_source_count;
  reg [5-1:0] _stream_conv2d_4_source_41_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_41_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_41_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_41_source_size;
  reg [32-1:0] _stream_conv2d_4_source_41_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_41_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_41_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_41_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_41_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_41_source_ram_raddr;
  reg _stream_conv2d_4_source_41_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_41_source_ram_rdata;
  reg _stream_conv2d_4_source_41_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_41_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_41_source_empty_data;
  reg _stream_conv2d_4_source_42_idle;
  reg [33-1:0] _stream_conv2d_4_source_42_source_count;
  reg [5-1:0] _stream_conv2d_4_source_42_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_42_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_42_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_42_source_size;
  reg [32-1:0] _stream_conv2d_4_source_42_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_42_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_42_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_42_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_42_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_42_source_ram_raddr;
  reg _stream_conv2d_4_source_42_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_42_source_ram_rdata;
  reg _stream_conv2d_4_source_42_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_42_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_42_source_empty_data;
  reg _stream_conv2d_4_source_43_idle;
  reg [33-1:0] _stream_conv2d_4_source_43_source_count;
  reg [5-1:0] _stream_conv2d_4_source_43_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_43_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_43_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_43_source_size;
  reg [32-1:0] _stream_conv2d_4_source_43_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_43_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_43_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_43_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_43_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_43_source_ram_raddr;
  reg _stream_conv2d_4_source_43_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_43_source_ram_rdata;
  reg _stream_conv2d_4_source_43_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_43_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_43_source_empty_data;
  reg _stream_conv2d_4_source_44_idle;
  reg [33-1:0] _stream_conv2d_4_source_44_source_count;
  reg [5-1:0] _stream_conv2d_4_source_44_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_44_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_44_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_44_source_size;
  reg [32-1:0] _stream_conv2d_4_source_44_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_44_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_44_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_44_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_44_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_44_source_ram_raddr;
  reg _stream_conv2d_4_source_44_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_44_source_ram_rdata;
  reg _stream_conv2d_4_source_44_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_44_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_44_source_empty_data;
  reg _stream_conv2d_4_source_45_idle;
  reg [33-1:0] _stream_conv2d_4_source_45_source_count;
  reg [5-1:0] _stream_conv2d_4_source_45_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_45_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_45_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_45_source_size;
  reg [32-1:0] _stream_conv2d_4_source_45_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_45_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_45_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_45_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_45_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_45_source_ram_raddr;
  reg _stream_conv2d_4_source_45_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_45_source_ram_rdata;
  reg _stream_conv2d_4_source_45_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_45_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_45_source_empty_data;
  reg _stream_conv2d_4_source_46_idle;
  reg [33-1:0] _stream_conv2d_4_source_46_source_count;
  reg [5-1:0] _stream_conv2d_4_source_46_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_46_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_46_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_46_source_size;
  reg [32-1:0] _stream_conv2d_4_source_46_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_46_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_46_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_46_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_46_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_46_source_ram_raddr;
  reg _stream_conv2d_4_source_46_source_ram_renable;
  wire [32-1:0] _stream_conv2d_4_source_46_source_ram_rdata;
  reg _stream_conv2d_4_source_46_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_4_source_46_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_4_source_46_source_empty_data;
  wire signed [16-1:0] mul_8_x_data;
  wire signed [16-1:0] mul_8_y_data;
  wire [5-1:0] mul_8_rshift_data;
  reg __mul_8_stream_ivalid_1;
  reg __mul_8_stream_ivalid_2;
  reg __mul_8_stream_ivalid_3;
  reg __mul_8_stream_ivalid_4;
  reg __mul_8_stream_ivalid_5;
  reg __mul_8_stream_ivalid_6;
  reg __mul_8_stream_ivalid_7;
  reg __mul_8_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_179;
  reg [5-1:0] _minus_data_181;
  reg [1-1:0] _greatereq_data_192;
  reg signed [16-1:0] __delay_data_1602__variable_176;
  reg signed [16-1:0] __delay_data_1605__variable_177;
  reg [5-1:0] __delay_data_1608__variable_178;
  reg signed [34-1:0] _sll_data_183;
  reg [1-1:0] __delay_data_1599_greaterthan_179;
  reg [1-1:0] __delay_data_1600_greatereq_192;
  reg signed [16-1:0] __delay_data_1603__delay_1602__variable_176;
  reg signed [16-1:0] __delay_data_1606__delay_1605__variable_177;
  reg [5-1:0] __delay_data_1609__delay_1608__variable_178;
  reg signed [32-1:0] _cond_data_189;
  reg [1-1:0] __delay_data_1601__delay_1600_greatereq_192;
  reg signed [16-1:0] __delay_data_1604__delay_1603__delay_1602__variable_176;
  reg signed [16-1:0] __delay_data_1607__delay_1606__delay_1605__variable_177;
  reg [5-1:0] __delay_data_1610__delay_1609__delay_1608__variable_178;
  wire signed [16-1:0] _uminus_data_191;
  assign _uminus_data_191 = -_cond_data_189;
  wire signed [16-1:0] _cond_data_194;
  assign _cond_data_194 = (__delay_data_1601__delay_1600_greatereq_192)? _cond_data_189 : _uminus_data_191;
  wire signed [32-1:0] __muladd_madd_odata_195;
  reg signed [32-1:0] __muladd_madd_odata_reg_195;
  wire signed [32-1:0] __muladd_data_195;
  assign __muladd_data_195 = __muladd_madd_odata_reg_195;
  wire __muladd_madd_update_195;
  assign __muladd_madd_update_195 = _mul_8_stream_oready;

  madd_0
  __muladd_madd_195
  (
    .CLK(CLK),
    .update(__muladd_madd_update_195),
    .a(__delay_data_1604__delay_1603__delay_1602__variable_176),
    .b(__delay_data_1607__delay_1606__delay_1605__variable_177),
    .c(_cond_data_194),
    .d(__muladd_madd_odata_195)
  );

  reg [5-1:0] __delay_data_1611__delay_1610__delay_1609____variable_178;
  reg [5-1:0] __delay_data_1612__delay_1611__delay_1610____variable_178;
  reg [5-1:0] __delay_data_1613__delay_1612__delay_1611____variable_178;
  reg [5-1:0] __delay_data_1614__delay_1613__delay_1612____variable_178;
  reg signed [32-1:0] _sra_data_196;
  wire signed [32-1:0] mul_8_z_data;
  assign mul_8_z_data = _sra_data_196;
  wire signed [16-1:0] mul_9_x_data;
  wire signed [16-1:0] mul_9_y_data;
  wire [5-1:0] mul_9_rshift_data;
  reg __mul_9_stream_ivalid_1;
  reg __mul_9_stream_ivalid_2;
  reg __mul_9_stream_ivalid_3;
  reg __mul_9_stream_ivalid_4;
  reg __mul_9_stream_ivalid_5;
  reg __mul_9_stream_ivalid_6;
  reg __mul_9_stream_ivalid_7;
  reg __mul_9_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_200;
  reg [5-1:0] _minus_data_202;
  reg [1-1:0] _greatereq_data_213;
  reg signed [16-1:0] __delay_data_1621__variable_197;
  reg signed [16-1:0] __delay_data_1624__variable_198;
  reg [5-1:0] __delay_data_1627__variable_199;
  reg signed [34-1:0] _sll_data_204;
  reg [1-1:0] __delay_data_1618_greaterthan_200;
  reg [1-1:0] __delay_data_1619_greatereq_213;
  reg signed [16-1:0] __delay_data_1622__delay_1621__variable_197;
  reg signed [16-1:0] __delay_data_1625__delay_1624__variable_198;
  reg [5-1:0] __delay_data_1628__delay_1627__variable_199;
  reg signed [32-1:0] _cond_data_210;
  reg [1-1:0] __delay_data_1620__delay_1619_greatereq_213;
  reg signed [16-1:0] __delay_data_1623__delay_1622__delay_1621__variable_197;
  reg signed [16-1:0] __delay_data_1626__delay_1625__delay_1624__variable_198;
  reg [5-1:0] __delay_data_1629__delay_1628__delay_1627__variable_199;
  wire signed [16-1:0] _uminus_data_212;
  assign _uminus_data_212 = -_cond_data_210;
  wire signed [16-1:0] _cond_data_215;
  assign _cond_data_215 = (__delay_data_1620__delay_1619_greatereq_213)? _cond_data_210 : _uminus_data_212;
  wire signed [32-1:0] __muladd_madd_odata_216;
  reg signed [32-1:0] __muladd_madd_odata_reg_216;
  wire signed [32-1:0] __muladd_data_216;
  assign __muladd_data_216 = __muladd_madd_odata_reg_216;
  wire __muladd_madd_update_216;
  assign __muladd_madd_update_216 = _mul_9_stream_oready;

  madd_1
  __muladd_madd_216
  (
    .CLK(CLK),
    .update(__muladd_madd_update_216),
    .a(__delay_data_1623__delay_1622__delay_1621__variable_197),
    .b(__delay_data_1626__delay_1625__delay_1624__variable_198),
    .c(_cond_data_215),
    .d(__muladd_madd_odata_216)
  );

  reg [5-1:0] __delay_data_1630__delay_1629__delay_1628____variable_199;
  reg [5-1:0] __delay_data_1631__delay_1630__delay_1629____variable_199;
  reg [5-1:0] __delay_data_1632__delay_1631__delay_1630____variable_199;
  reg [5-1:0] __delay_data_1633__delay_1632__delay_1631____variable_199;
  reg signed [32-1:0] _sra_data_217;
  wire signed [32-1:0] mul_9_z_data;
  assign mul_9_z_data = _sra_data_217;
  wire signed [16-1:0] mul_10_x_data;
  wire signed [16-1:0] mul_10_y_data;
  wire [5-1:0] mul_10_rshift_data;
  reg __mul_10_stream_ivalid_1;
  reg __mul_10_stream_ivalid_2;
  reg __mul_10_stream_ivalid_3;
  reg __mul_10_stream_ivalid_4;
  reg __mul_10_stream_ivalid_5;
  reg __mul_10_stream_ivalid_6;
  reg __mul_10_stream_ivalid_7;
  reg __mul_10_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_221;
  reg [5-1:0] _minus_data_223;
  reg [1-1:0] _greatereq_data_234;
  reg signed [16-1:0] __delay_data_1640__variable_218;
  reg signed [16-1:0] __delay_data_1643__variable_219;
  reg [5-1:0] __delay_data_1646__variable_220;
  reg signed [34-1:0] _sll_data_225;
  reg [1-1:0] __delay_data_1637_greaterthan_221;
  reg [1-1:0] __delay_data_1638_greatereq_234;
  reg signed [16-1:0] __delay_data_1641__delay_1640__variable_218;
  reg signed [16-1:0] __delay_data_1644__delay_1643__variable_219;
  reg [5-1:0] __delay_data_1647__delay_1646__variable_220;
  reg signed [32-1:0] _cond_data_231;
  reg [1-1:0] __delay_data_1639__delay_1638_greatereq_234;
  reg signed [16-1:0] __delay_data_1642__delay_1641__delay_1640__variable_218;
  reg signed [16-1:0] __delay_data_1645__delay_1644__delay_1643__variable_219;
  reg [5-1:0] __delay_data_1648__delay_1647__delay_1646__variable_220;
  wire signed [16-1:0] _uminus_data_233;
  assign _uminus_data_233 = -_cond_data_231;
  wire signed [16-1:0] _cond_data_236;
  assign _cond_data_236 = (__delay_data_1639__delay_1638_greatereq_234)? _cond_data_231 : _uminus_data_233;
  wire signed [32-1:0] __muladd_madd_odata_237;
  reg signed [32-1:0] __muladd_madd_odata_reg_237;
  wire signed [32-1:0] __muladd_data_237;
  assign __muladd_data_237 = __muladd_madd_odata_reg_237;
  wire __muladd_madd_update_237;
  assign __muladd_madd_update_237 = _mul_10_stream_oready;

  madd_2
  __muladd_madd_237
  (
    .CLK(CLK),
    .update(__muladd_madd_update_237),
    .a(__delay_data_1642__delay_1641__delay_1640__variable_218),
    .b(__delay_data_1645__delay_1644__delay_1643__variable_219),
    .c(_cond_data_236),
    .d(__muladd_madd_odata_237)
  );

  reg [5-1:0] __delay_data_1649__delay_1648__delay_1647____variable_220;
  reg [5-1:0] __delay_data_1650__delay_1649__delay_1648____variable_220;
  reg [5-1:0] __delay_data_1651__delay_1650__delay_1649____variable_220;
  reg [5-1:0] __delay_data_1652__delay_1651__delay_1650____variable_220;
  reg signed [32-1:0] _sra_data_238;
  wire signed [32-1:0] mul_10_z_data;
  assign mul_10_z_data = _sra_data_238;
  wire signed [16-1:0] mul_11_x_data;
  wire signed [16-1:0] mul_11_y_data;
  wire [5-1:0] mul_11_rshift_data;
  reg __mul_11_stream_ivalid_1;
  reg __mul_11_stream_ivalid_2;
  reg __mul_11_stream_ivalid_3;
  reg __mul_11_stream_ivalid_4;
  reg __mul_11_stream_ivalid_5;
  reg __mul_11_stream_ivalid_6;
  reg __mul_11_stream_ivalid_7;
  reg __mul_11_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_242;
  reg [5-1:0] _minus_data_244;
  reg [1-1:0] _greatereq_data_255;
  reg signed [16-1:0] __delay_data_1659__variable_239;
  reg signed [16-1:0] __delay_data_1662__variable_240;
  reg [5-1:0] __delay_data_1665__variable_241;
  reg signed [34-1:0] _sll_data_246;
  reg [1-1:0] __delay_data_1656_greaterthan_242;
  reg [1-1:0] __delay_data_1657_greatereq_255;
  reg signed [16-1:0] __delay_data_1660__delay_1659__variable_239;
  reg signed [16-1:0] __delay_data_1663__delay_1662__variable_240;
  reg [5-1:0] __delay_data_1666__delay_1665__variable_241;
  reg signed [32-1:0] _cond_data_252;
  reg [1-1:0] __delay_data_1658__delay_1657_greatereq_255;
  reg signed [16-1:0] __delay_data_1661__delay_1660__delay_1659__variable_239;
  reg signed [16-1:0] __delay_data_1664__delay_1663__delay_1662__variable_240;
  reg [5-1:0] __delay_data_1667__delay_1666__delay_1665__variable_241;
  wire signed [16-1:0] _uminus_data_254;
  assign _uminus_data_254 = -_cond_data_252;
  wire signed [16-1:0] _cond_data_257;
  assign _cond_data_257 = (__delay_data_1658__delay_1657_greatereq_255)? _cond_data_252 : _uminus_data_254;
  wire signed [32-1:0] __muladd_madd_odata_258;
  reg signed [32-1:0] __muladd_madd_odata_reg_258;
  wire signed [32-1:0] __muladd_data_258;
  assign __muladd_data_258 = __muladd_madd_odata_reg_258;
  wire __muladd_madd_update_258;
  assign __muladd_madd_update_258 = _mul_11_stream_oready;

  madd_3
  __muladd_madd_258
  (
    .CLK(CLK),
    .update(__muladd_madd_update_258),
    .a(__delay_data_1661__delay_1660__delay_1659__variable_239),
    .b(__delay_data_1664__delay_1663__delay_1662__variable_240),
    .c(_cond_data_257),
    .d(__muladd_madd_odata_258)
  );

  reg [5-1:0] __delay_data_1668__delay_1667__delay_1666____variable_241;
  reg [5-1:0] __delay_data_1669__delay_1668__delay_1667____variable_241;
  reg [5-1:0] __delay_data_1670__delay_1669__delay_1668____variable_241;
  reg [5-1:0] __delay_data_1671__delay_1670__delay_1669____variable_241;
  reg signed [32-1:0] _sra_data_259;
  wire signed [32-1:0] mul_11_z_data;
  assign mul_11_z_data = _sra_data_259;
  wire signed [16-1:0] mul_12_x_data;
  wire signed [16-1:0] mul_12_y_data;
  wire [5-1:0] mul_12_rshift_data;
  reg __mul_12_stream_ivalid_1;
  reg __mul_12_stream_ivalid_2;
  reg __mul_12_stream_ivalid_3;
  reg __mul_12_stream_ivalid_4;
  reg __mul_12_stream_ivalid_5;
  reg __mul_12_stream_ivalid_6;
  reg __mul_12_stream_ivalid_7;
  reg __mul_12_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_263;
  reg [5-1:0] _minus_data_265;
  reg [1-1:0] _greatereq_data_276;
  reg signed [16-1:0] __delay_data_1678__variable_260;
  reg signed [16-1:0] __delay_data_1681__variable_261;
  reg [5-1:0] __delay_data_1684__variable_262;
  reg signed [34-1:0] _sll_data_267;
  reg [1-1:0] __delay_data_1675_greaterthan_263;
  reg [1-1:0] __delay_data_1676_greatereq_276;
  reg signed [16-1:0] __delay_data_1679__delay_1678__variable_260;
  reg signed [16-1:0] __delay_data_1682__delay_1681__variable_261;
  reg [5-1:0] __delay_data_1685__delay_1684__variable_262;
  reg signed [32-1:0] _cond_data_273;
  reg [1-1:0] __delay_data_1677__delay_1676_greatereq_276;
  reg signed [16-1:0] __delay_data_1680__delay_1679__delay_1678__variable_260;
  reg signed [16-1:0] __delay_data_1683__delay_1682__delay_1681__variable_261;
  reg [5-1:0] __delay_data_1686__delay_1685__delay_1684__variable_262;
  wire signed [16-1:0] _uminus_data_275;
  assign _uminus_data_275 = -_cond_data_273;
  wire signed [16-1:0] _cond_data_278;
  assign _cond_data_278 = (__delay_data_1677__delay_1676_greatereq_276)? _cond_data_273 : _uminus_data_275;
  wire signed [32-1:0] __muladd_madd_odata_279;
  reg signed [32-1:0] __muladd_madd_odata_reg_279;
  wire signed [32-1:0] __muladd_data_279;
  assign __muladd_data_279 = __muladd_madd_odata_reg_279;
  wire __muladd_madd_update_279;
  assign __muladd_madd_update_279 = _mul_12_stream_oready;

  madd_4
  __muladd_madd_279
  (
    .CLK(CLK),
    .update(__muladd_madd_update_279),
    .a(__delay_data_1680__delay_1679__delay_1678__variable_260),
    .b(__delay_data_1683__delay_1682__delay_1681__variable_261),
    .c(_cond_data_278),
    .d(__muladd_madd_odata_279)
  );

  reg [5-1:0] __delay_data_1687__delay_1686__delay_1685____variable_262;
  reg [5-1:0] __delay_data_1688__delay_1687__delay_1686____variable_262;
  reg [5-1:0] __delay_data_1689__delay_1688__delay_1687____variable_262;
  reg [5-1:0] __delay_data_1690__delay_1689__delay_1688____variable_262;
  reg signed [32-1:0] _sra_data_280;
  wire signed [32-1:0] mul_12_z_data;
  assign mul_12_z_data = _sra_data_280;
  wire signed [16-1:0] mul_13_x_data;
  wire signed [16-1:0] mul_13_y_data;
  wire [5-1:0] mul_13_rshift_data;
  reg __mul_13_stream_ivalid_1;
  reg __mul_13_stream_ivalid_2;
  reg __mul_13_stream_ivalid_3;
  reg __mul_13_stream_ivalid_4;
  reg __mul_13_stream_ivalid_5;
  reg __mul_13_stream_ivalid_6;
  reg __mul_13_stream_ivalid_7;
  reg __mul_13_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_284;
  reg [5-1:0] _minus_data_286;
  reg [1-1:0] _greatereq_data_297;
  reg signed [16-1:0] __delay_data_1697__variable_281;
  reg signed [16-1:0] __delay_data_1700__variable_282;
  reg [5-1:0] __delay_data_1703__variable_283;
  reg signed [34-1:0] _sll_data_288;
  reg [1-1:0] __delay_data_1694_greaterthan_284;
  reg [1-1:0] __delay_data_1695_greatereq_297;
  reg signed [16-1:0] __delay_data_1698__delay_1697__variable_281;
  reg signed [16-1:0] __delay_data_1701__delay_1700__variable_282;
  reg [5-1:0] __delay_data_1704__delay_1703__variable_283;
  reg signed [32-1:0] _cond_data_294;
  reg [1-1:0] __delay_data_1696__delay_1695_greatereq_297;
  reg signed [16-1:0] __delay_data_1699__delay_1698__delay_1697__variable_281;
  reg signed [16-1:0] __delay_data_1702__delay_1701__delay_1700__variable_282;
  reg [5-1:0] __delay_data_1705__delay_1704__delay_1703__variable_283;
  wire signed [16-1:0] _uminus_data_296;
  assign _uminus_data_296 = -_cond_data_294;
  wire signed [16-1:0] _cond_data_299;
  assign _cond_data_299 = (__delay_data_1696__delay_1695_greatereq_297)? _cond_data_294 : _uminus_data_296;
  wire signed [32-1:0] __muladd_madd_odata_300;
  reg signed [32-1:0] __muladd_madd_odata_reg_300;
  wire signed [32-1:0] __muladd_data_300;
  assign __muladd_data_300 = __muladd_madd_odata_reg_300;
  wire __muladd_madd_update_300;
  assign __muladd_madd_update_300 = _mul_13_stream_oready;

  madd_5
  __muladd_madd_300
  (
    .CLK(CLK),
    .update(__muladd_madd_update_300),
    .a(__delay_data_1699__delay_1698__delay_1697__variable_281),
    .b(__delay_data_1702__delay_1701__delay_1700__variable_282),
    .c(_cond_data_299),
    .d(__muladd_madd_odata_300)
  );

  reg [5-1:0] __delay_data_1706__delay_1705__delay_1704____variable_283;
  reg [5-1:0] __delay_data_1707__delay_1706__delay_1705____variable_283;
  reg [5-1:0] __delay_data_1708__delay_1707__delay_1706____variable_283;
  reg [5-1:0] __delay_data_1709__delay_1708__delay_1707____variable_283;
  reg signed [32-1:0] _sra_data_301;
  wire signed [32-1:0] mul_13_z_data;
  assign mul_13_z_data = _sra_data_301;
  wire signed [16-1:0] mul_14_x_data;
  wire signed [16-1:0] mul_14_y_data;
  wire [5-1:0] mul_14_rshift_data;
  reg __mul_14_stream_ivalid_1;
  reg __mul_14_stream_ivalid_2;
  reg __mul_14_stream_ivalid_3;
  reg __mul_14_stream_ivalid_4;
  reg __mul_14_stream_ivalid_5;
  reg __mul_14_stream_ivalid_6;
  reg __mul_14_stream_ivalid_7;
  reg __mul_14_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_305;
  reg [5-1:0] _minus_data_307;
  reg [1-1:0] _greatereq_data_318;
  reg signed [16-1:0] __delay_data_1716__variable_302;
  reg signed [16-1:0] __delay_data_1719__variable_303;
  reg [5-1:0] __delay_data_1722__variable_304;
  reg signed [34-1:0] _sll_data_309;
  reg [1-1:0] __delay_data_1713_greaterthan_305;
  reg [1-1:0] __delay_data_1714_greatereq_318;
  reg signed [16-1:0] __delay_data_1717__delay_1716__variable_302;
  reg signed [16-1:0] __delay_data_1720__delay_1719__variable_303;
  reg [5-1:0] __delay_data_1723__delay_1722__variable_304;
  reg signed [32-1:0] _cond_data_315;
  reg [1-1:0] __delay_data_1715__delay_1714_greatereq_318;
  reg signed [16-1:0] __delay_data_1718__delay_1717__delay_1716__variable_302;
  reg signed [16-1:0] __delay_data_1721__delay_1720__delay_1719__variable_303;
  reg [5-1:0] __delay_data_1724__delay_1723__delay_1722__variable_304;
  wire signed [16-1:0] _uminus_data_317;
  assign _uminus_data_317 = -_cond_data_315;
  wire signed [16-1:0] _cond_data_320;
  assign _cond_data_320 = (__delay_data_1715__delay_1714_greatereq_318)? _cond_data_315 : _uminus_data_317;
  wire signed [32-1:0] __muladd_madd_odata_321;
  reg signed [32-1:0] __muladd_madd_odata_reg_321;
  wire signed [32-1:0] __muladd_data_321;
  assign __muladd_data_321 = __muladd_madd_odata_reg_321;
  wire __muladd_madd_update_321;
  assign __muladd_madd_update_321 = _mul_14_stream_oready;

  madd_6
  __muladd_madd_321
  (
    .CLK(CLK),
    .update(__muladd_madd_update_321),
    .a(__delay_data_1718__delay_1717__delay_1716__variable_302),
    .b(__delay_data_1721__delay_1720__delay_1719__variable_303),
    .c(_cond_data_320),
    .d(__muladd_madd_odata_321)
  );

  reg [5-1:0] __delay_data_1725__delay_1724__delay_1723____variable_304;
  reg [5-1:0] __delay_data_1726__delay_1725__delay_1724____variable_304;
  reg [5-1:0] __delay_data_1727__delay_1726__delay_1725____variable_304;
  reg [5-1:0] __delay_data_1728__delay_1727__delay_1726____variable_304;
  reg signed [32-1:0] _sra_data_322;
  wire signed [32-1:0] mul_14_z_data;
  assign mul_14_z_data = _sra_data_322;
  wire signed [16-1:0] mul_15_x_data;
  wire signed [16-1:0] mul_15_y_data;
  wire [5-1:0] mul_15_rshift_data;
  reg __mul_15_stream_ivalid_1;
  reg __mul_15_stream_ivalid_2;
  reg __mul_15_stream_ivalid_3;
  reg __mul_15_stream_ivalid_4;
  reg __mul_15_stream_ivalid_5;
  reg __mul_15_stream_ivalid_6;
  reg __mul_15_stream_ivalid_7;
  reg __mul_15_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_326;
  reg [5-1:0] _minus_data_328;
  reg [1-1:0] _greatereq_data_339;
  reg signed [16-1:0] __delay_data_1735__variable_323;
  reg signed [16-1:0] __delay_data_1738__variable_324;
  reg [5-1:0] __delay_data_1741__variable_325;
  reg signed [34-1:0] _sll_data_330;
  reg [1-1:0] __delay_data_1732_greaterthan_326;
  reg [1-1:0] __delay_data_1733_greatereq_339;
  reg signed [16-1:0] __delay_data_1736__delay_1735__variable_323;
  reg signed [16-1:0] __delay_data_1739__delay_1738__variable_324;
  reg [5-1:0] __delay_data_1742__delay_1741__variable_325;
  reg signed [32-1:0] _cond_data_336;
  reg [1-1:0] __delay_data_1734__delay_1733_greatereq_339;
  reg signed [16-1:0] __delay_data_1737__delay_1736__delay_1735__variable_323;
  reg signed [16-1:0] __delay_data_1740__delay_1739__delay_1738__variable_324;
  reg [5-1:0] __delay_data_1743__delay_1742__delay_1741__variable_325;
  wire signed [16-1:0] _uminus_data_338;
  assign _uminus_data_338 = -_cond_data_336;
  wire signed [16-1:0] _cond_data_341;
  assign _cond_data_341 = (__delay_data_1734__delay_1733_greatereq_339)? _cond_data_336 : _uminus_data_338;
  wire signed [32-1:0] __muladd_madd_odata_342;
  reg signed [32-1:0] __muladd_madd_odata_reg_342;
  wire signed [32-1:0] __muladd_data_342;
  assign __muladd_data_342 = __muladd_madd_odata_reg_342;
  wire __muladd_madd_update_342;
  assign __muladd_madd_update_342 = _mul_15_stream_oready;

  madd_7
  __muladd_madd_342
  (
    .CLK(CLK),
    .update(__muladd_madd_update_342),
    .a(__delay_data_1737__delay_1736__delay_1735__variable_323),
    .b(__delay_data_1740__delay_1739__delay_1738__variable_324),
    .c(_cond_data_341),
    .d(__muladd_madd_odata_342)
  );

  reg [5-1:0] __delay_data_1744__delay_1743__delay_1742____variable_325;
  reg [5-1:0] __delay_data_1745__delay_1744__delay_1743____variable_325;
  reg [5-1:0] __delay_data_1746__delay_1745__delay_1744____variable_325;
  reg [5-1:0] __delay_data_1747__delay_1746__delay_1745____variable_325;
  reg signed [32-1:0] _sra_data_343;
  wire signed [32-1:0] mul_15_z_data;
  assign mul_15_z_data = _sra_data_343;
  wire signed [16-1:0] mul_16_x_data;
  wire signed [16-1:0] mul_16_y_data;
  wire [5-1:0] mul_16_rshift_data;
  reg __mul_16_stream_ivalid_1;
  reg __mul_16_stream_ivalid_2;
  reg __mul_16_stream_ivalid_3;
  reg __mul_16_stream_ivalid_4;
  reg __mul_16_stream_ivalid_5;
  reg __mul_16_stream_ivalid_6;
  reg __mul_16_stream_ivalid_7;
  reg __mul_16_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_347;
  reg [5-1:0] _minus_data_349;
  reg [1-1:0] _greatereq_data_360;
  reg signed [16-1:0] __delay_data_1754__variable_344;
  reg signed [16-1:0] __delay_data_1757__variable_345;
  reg [5-1:0] __delay_data_1760__variable_346;
  reg signed [34-1:0] _sll_data_351;
  reg [1-1:0] __delay_data_1751_greaterthan_347;
  reg [1-1:0] __delay_data_1752_greatereq_360;
  reg signed [16-1:0] __delay_data_1755__delay_1754__variable_344;
  reg signed [16-1:0] __delay_data_1758__delay_1757__variable_345;
  reg [5-1:0] __delay_data_1761__delay_1760__variable_346;
  reg signed [32-1:0] _cond_data_357;
  reg [1-1:0] __delay_data_1753__delay_1752_greatereq_360;
  reg signed [16-1:0] __delay_data_1756__delay_1755__delay_1754__variable_344;
  reg signed [16-1:0] __delay_data_1759__delay_1758__delay_1757__variable_345;
  reg [5-1:0] __delay_data_1762__delay_1761__delay_1760__variable_346;
  wire signed [16-1:0] _uminus_data_359;
  assign _uminus_data_359 = -_cond_data_357;
  wire signed [16-1:0] _cond_data_362;
  assign _cond_data_362 = (__delay_data_1753__delay_1752_greatereq_360)? _cond_data_357 : _uminus_data_359;
  wire signed [32-1:0] __muladd_madd_odata_363;
  reg signed [32-1:0] __muladd_madd_odata_reg_363;
  wire signed [32-1:0] __muladd_data_363;
  assign __muladd_data_363 = __muladd_madd_odata_reg_363;
  wire __muladd_madd_update_363;
  assign __muladd_madd_update_363 = _mul_16_stream_oready;

  madd_8
  __muladd_madd_363
  (
    .CLK(CLK),
    .update(__muladd_madd_update_363),
    .a(__delay_data_1756__delay_1755__delay_1754__variable_344),
    .b(__delay_data_1759__delay_1758__delay_1757__variable_345),
    .c(_cond_data_362),
    .d(__muladd_madd_odata_363)
  );

  reg [5-1:0] __delay_data_1763__delay_1762__delay_1761____variable_346;
  reg [5-1:0] __delay_data_1764__delay_1763__delay_1762____variable_346;
  reg [5-1:0] __delay_data_1765__delay_1764__delay_1763____variable_346;
  reg [5-1:0] __delay_data_1766__delay_1765__delay_1764____variable_346;
  reg signed [32-1:0] _sra_data_364;
  wire signed [32-1:0] mul_16_z_data;
  assign mul_16_z_data = _sra_data_364;
  wire signed [16-1:0] mul_17_x_data;
  wire signed [16-1:0] mul_17_y_data;
  wire [5-1:0] mul_17_rshift_data;
  reg __mul_17_stream_ivalid_1;
  reg __mul_17_stream_ivalid_2;
  reg __mul_17_stream_ivalid_3;
  reg __mul_17_stream_ivalid_4;
  reg __mul_17_stream_ivalid_5;
  reg __mul_17_stream_ivalid_6;
  reg __mul_17_stream_ivalid_7;
  reg __mul_17_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_368;
  reg [5-1:0] _minus_data_370;
  reg [1-1:0] _greatereq_data_381;
  reg signed [16-1:0] __delay_data_1791__variable_365;
  reg signed [16-1:0] __delay_data_1794__variable_366;
  reg [5-1:0] __delay_data_1797__variable_367;
  reg signed [34-1:0] _sll_data_372;
  reg [1-1:0] __delay_data_1788_greaterthan_368;
  reg [1-1:0] __delay_data_1789_greatereq_381;
  reg signed [16-1:0] __delay_data_1792__delay_1791__variable_365;
  reg signed [16-1:0] __delay_data_1795__delay_1794__variable_366;
  reg [5-1:0] __delay_data_1798__delay_1797__variable_367;
  reg signed [32-1:0] _cond_data_378;
  reg [1-1:0] __delay_data_1790__delay_1789_greatereq_381;
  reg signed [16-1:0] __delay_data_1793__delay_1792__delay_1791__variable_365;
  reg signed [16-1:0] __delay_data_1796__delay_1795__delay_1794__variable_366;
  reg [5-1:0] __delay_data_1799__delay_1798__delay_1797__variable_367;
  wire signed [16-1:0] _uminus_data_380;
  assign _uminus_data_380 = -_cond_data_378;
  wire signed [16-1:0] _cond_data_383;
  assign _cond_data_383 = (__delay_data_1790__delay_1789_greatereq_381)? _cond_data_378 : _uminus_data_380;
  wire signed [32-1:0] __muladd_madd_odata_384;
  reg signed [32-1:0] __muladd_madd_odata_reg_384;
  wire signed [32-1:0] __muladd_data_384;
  assign __muladd_data_384 = __muladd_madd_odata_reg_384;
  wire __muladd_madd_update_384;
  assign __muladd_madd_update_384 = _mul_17_stream_oready;

  madd_9
  __muladd_madd_384
  (
    .CLK(CLK),
    .update(__muladd_madd_update_384),
    .a(__delay_data_1793__delay_1792__delay_1791__variable_365),
    .b(__delay_data_1796__delay_1795__delay_1794__variable_366),
    .c(_cond_data_383),
    .d(__muladd_madd_odata_384)
  );

  reg [5-1:0] __delay_data_1800__delay_1799__delay_1798____variable_367;
  reg [5-1:0] __delay_data_1801__delay_1800__delay_1799____variable_367;
  reg [5-1:0] __delay_data_1802__delay_1801__delay_1800____variable_367;
  reg [5-1:0] __delay_data_1803__delay_1802__delay_1801____variable_367;
  reg signed [32-1:0] _sra_data_385;
  wire signed [32-1:0] mul_17_z_data;
  assign mul_17_z_data = _sra_data_385;
  wire signed [16-1:0] mul_18_x_data;
  wire signed [16-1:0] mul_18_y_data;
  wire [5-1:0] mul_18_rshift_data;
  reg __mul_18_stream_ivalid_1;
  reg __mul_18_stream_ivalid_2;
  reg __mul_18_stream_ivalid_3;
  reg __mul_18_stream_ivalid_4;
  reg __mul_18_stream_ivalid_5;
  reg __mul_18_stream_ivalid_6;
  reg __mul_18_stream_ivalid_7;
  reg __mul_18_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_389;
  reg [5-1:0] _minus_data_391;
  reg [1-1:0] _greatereq_data_402;
  reg signed [16-1:0] __delay_data_1810__variable_386;
  reg signed [16-1:0] __delay_data_1813__variable_387;
  reg [5-1:0] __delay_data_1816__variable_388;
  reg signed [34-1:0] _sll_data_393;
  reg [1-1:0] __delay_data_1807_greaterthan_389;
  reg [1-1:0] __delay_data_1808_greatereq_402;
  reg signed [16-1:0] __delay_data_1811__delay_1810__variable_386;
  reg signed [16-1:0] __delay_data_1814__delay_1813__variable_387;
  reg [5-1:0] __delay_data_1817__delay_1816__variable_388;
  reg signed [32-1:0] _cond_data_399;
  reg [1-1:0] __delay_data_1809__delay_1808_greatereq_402;
  reg signed [16-1:0] __delay_data_1812__delay_1811__delay_1810__variable_386;
  reg signed [16-1:0] __delay_data_1815__delay_1814__delay_1813__variable_387;
  reg [5-1:0] __delay_data_1818__delay_1817__delay_1816__variable_388;
  wire signed [16-1:0] _uminus_data_401;
  assign _uminus_data_401 = -_cond_data_399;
  wire signed [16-1:0] _cond_data_404;
  assign _cond_data_404 = (__delay_data_1809__delay_1808_greatereq_402)? _cond_data_399 : _uminus_data_401;
  wire signed [32-1:0] __muladd_madd_odata_405;
  reg signed [32-1:0] __muladd_madd_odata_reg_405;
  wire signed [32-1:0] __muladd_data_405;
  assign __muladd_data_405 = __muladd_madd_odata_reg_405;
  wire __muladd_madd_update_405;
  assign __muladd_madd_update_405 = _mul_18_stream_oready;

  madd_10
  __muladd_madd_405
  (
    .CLK(CLK),
    .update(__muladd_madd_update_405),
    .a(__delay_data_1812__delay_1811__delay_1810__variable_386),
    .b(__delay_data_1815__delay_1814__delay_1813__variable_387),
    .c(_cond_data_404),
    .d(__muladd_madd_odata_405)
  );

  reg [5-1:0] __delay_data_1819__delay_1818__delay_1817____variable_388;
  reg [5-1:0] __delay_data_1820__delay_1819__delay_1818____variable_388;
  reg [5-1:0] __delay_data_1821__delay_1820__delay_1819____variable_388;
  reg [5-1:0] __delay_data_1822__delay_1821__delay_1820____variable_388;
  reg signed [32-1:0] _sra_data_406;
  wire signed [32-1:0] mul_18_z_data;
  assign mul_18_z_data = _sra_data_406;
  wire signed [16-1:0] mul_19_x_data;
  wire signed [16-1:0] mul_19_y_data;
  wire [5-1:0] mul_19_rshift_data;
  reg __mul_19_stream_ivalid_1;
  reg __mul_19_stream_ivalid_2;
  reg __mul_19_stream_ivalid_3;
  reg __mul_19_stream_ivalid_4;
  reg __mul_19_stream_ivalid_5;
  reg __mul_19_stream_ivalid_6;
  reg __mul_19_stream_ivalid_7;
  reg __mul_19_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_410;
  reg [5-1:0] _minus_data_412;
  reg [1-1:0] _greatereq_data_423;
  reg signed [16-1:0] __delay_data_1829__variable_407;
  reg signed [16-1:0] __delay_data_1832__variable_408;
  reg [5-1:0] __delay_data_1835__variable_409;
  reg signed [34-1:0] _sll_data_414;
  reg [1-1:0] __delay_data_1826_greaterthan_410;
  reg [1-1:0] __delay_data_1827_greatereq_423;
  reg signed [16-1:0] __delay_data_1830__delay_1829__variable_407;
  reg signed [16-1:0] __delay_data_1833__delay_1832__variable_408;
  reg [5-1:0] __delay_data_1836__delay_1835__variable_409;
  reg signed [32-1:0] _cond_data_420;
  reg [1-1:0] __delay_data_1828__delay_1827_greatereq_423;
  reg signed [16-1:0] __delay_data_1831__delay_1830__delay_1829__variable_407;
  reg signed [16-1:0] __delay_data_1834__delay_1833__delay_1832__variable_408;
  reg [5-1:0] __delay_data_1837__delay_1836__delay_1835__variable_409;
  wire signed [16-1:0] _uminus_data_422;
  assign _uminus_data_422 = -_cond_data_420;
  wire signed [16-1:0] _cond_data_425;
  assign _cond_data_425 = (__delay_data_1828__delay_1827_greatereq_423)? _cond_data_420 : _uminus_data_422;
  wire signed [32-1:0] __muladd_madd_odata_426;
  reg signed [32-1:0] __muladd_madd_odata_reg_426;
  wire signed [32-1:0] __muladd_data_426;
  assign __muladd_data_426 = __muladd_madd_odata_reg_426;
  wire __muladd_madd_update_426;
  assign __muladd_madd_update_426 = _mul_19_stream_oready;

  madd_11
  __muladd_madd_426
  (
    .CLK(CLK),
    .update(__muladd_madd_update_426),
    .a(__delay_data_1831__delay_1830__delay_1829__variable_407),
    .b(__delay_data_1834__delay_1833__delay_1832__variable_408),
    .c(_cond_data_425),
    .d(__muladd_madd_odata_426)
  );

  reg [5-1:0] __delay_data_1838__delay_1837__delay_1836____variable_409;
  reg [5-1:0] __delay_data_1839__delay_1838__delay_1837____variable_409;
  reg [5-1:0] __delay_data_1840__delay_1839__delay_1838____variable_409;
  reg [5-1:0] __delay_data_1841__delay_1840__delay_1839____variable_409;
  reg signed [32-1:0] _sra_data_427;
  wire signed [32-1:0] mul_19_z_data;
  assign mul_19_z_data = _sra_data_427;
  wire signed [16-1:0] mul_20_x_data;
  wire signed [16-1:0] mul_20_y_data;
  wire [5-1:0] mul_20_rshift_data;
  reg __mul_20_stream_ivalid_1;
  reg __mul_20_stream_ivalid_2;
  reg __mul_20_stream_ivalid_3;
  reg __mul_20_stream_ivalid_4;
  reg __mul_20_stream_ivalid_5;
  reg __mul_20_stream_ivalid_6;
  reg __mul_20_stream_ivalid_7;
  reg __mul_20_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_431;
  reg [5-1:0] _minus_data_433;
  reg [1-1:0] _greatereq_data_444;
  reg signed [16-1:0] __delay_data_1848__variable_428;
  reg signed [16-1:0] __delay_data_1851__variable_429;
  reg [5-1:0] __delay_data_1854__variable_430;
  reg signed [34-1:0] _sll_data_435;
  reg [1-1:0] __delay_data_1845_greaterthan_431;
  reg [1-1:0] __delay_data_1846_greatereq_444;
  reg signed [16-1:0] __delay_data_1849__delay_1848__variable_428;
  reg signed [16-1:0] __delay_data_1852__delay_1851__variable_429;
  reg [5-1:0] __delay_data_1855__delay_1854__variable_430;
  reg signed [32-1:0] _cond_data_441;
  reg [1-1:0] __delay_data_1847__delay_1846_greatereq_444;
  reg signed [16-1:0] __delay_data_1850__delay_1849__delay_1848__variable_428;
  reg signed [16-1:0] __delay_data_1853__delay_1852__delay_1851__variable_429;
  reg [5-1:0] __delay_data_1856__delay_1855__delay_1854__variable_430;
  wire signed [16-1:0] _uminus_data_443;
  assign _uminus_data_443 = -_cond_data_441;
  wire signed [16-1:0] _cond_data_446;
  assign _cond_data_446 = (__delay_data_1847__delay_1846_greatereq_444)? _cond_data_441 : _uminus_data_443;
  wire signed [32-1:0] __muladd_madd_odata_447;
  reg signed [32-1:0] __muladd_madd_odata_reg_447;
  wire signed [32-1:0] __muladd_data_447;
  assign __muladd_data_447 = __muladd_madd_odata_reg_447;
  wire __muladd_madd_update_447;
  assign __muladd_madd_update_447 = _mul_20_stream_oready;

  madd_12
  __muladd_madd_447
  (
    .CLK(CLK),
    .update(__muladd_madd_update_447),
    .a(__delay_data_1850__delay_1849__delay_1848__variable_428),
    .b(__delay_data_1853__delay_1852__delay_1851__variable_429),
    .c(_cond_data_446),
    .d(__muladd_madd_odata_447)
  );

  reg [5-1:0] __delay_data_1857__delay_1856__delay_1855____variable_430;
  reg [5-1:0] __delay_data_1858__delay_1857__delay_1856____variable_430;
  reg [5-1:0] __delay_data_1859__delay_1858__delay_1857____variable_430;
  reg [5-1:0] __delay_data_1860__delay_1859__delay_1858____variable_430;
  reg signed [32-1:0] _sra_data_448;
  wire signed [32-1:0] mul_20_z_data;
  assign mul_20_z_data = _sra_data_448;
  wire signed [16-1:0] mul_21_x_data;
  wire signed [16-1:0] mul_21_y_data;
  wire [5-1:0] mul_21_rshift_data;
  reg __mul_21_stream_ivalid_1;
  reg __mul_21_stream_ivalid_2;
  reg __mul_21_stream_ivalid_3;
  reg __mul_21_stream_ivalid_4;
  reg __mul_21_stream_ivalid_5;
  reg __mul_21_stream_ivalid_6;
  reg __mul_21_stream_ivalid_7;
  reg __mul_21_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_452;
  reg [5-1:0] _minus_data_454;
  reg [1-1:0] _greatereq_data_465;
  reg signed [16-1:0] __delay_data_1867__variable_449;
  reg signed [16-1:0] __delay_data_1870__variable_450;
  reg [5-1:0] __delay_data_1873__variable_451;
  reg signed [34-1:0] _sll_data_456;
  reg [1-1:0] __delay_data_1864_greaterthan_452;
  reg [1-1:0] __delay_data_1865_greatereq_465;
  reg signed [16-1:0] __delay_data_1868__delay_1867__variable_449;
  reg signed [16-1:0] __delay_data_1871__delay_1870__variable_450;
  reg [5-1:0] __delay_data_1874__delay_1873__variable_451;
  reg signed [32-1:0] _cond_data_462;
  reg [1-1:0] __delay_data_1866__delay_1865_greatereq_465;
  reg signed [16-1:0] __delay_data_1869__delay_1868__delay_1867__variable_449;
  reg signed [16-1:0] __delay_data_1872__delay_1871__delay_1870__variable_450;
  reg [5-1:0] __delay_data_1875__delay_1874__delay_1873__variable_451;
  wire signed [16-1:0] _uminus_data_464;
  assign _uminus_data_464 = -_cond_data_462;
  wire signed [16-1:0] _cond_data_467;
  assign _cond_data_467 = (__delay_data_1866__delay_1865_greatereq_465)? _cond_data_462 : _uminus_data_464;
  wire signed [32-1:0] __muladd_madd_odata_468;
  reg signed [32-1:0] __muladd_madd_odata_reg_468;
  wire signed [32-1:0] __muladd_data_468;
  assign __muladd_data_468 = __muladd_madd_odata_reg_468;
  wire __muladd_madd_update_468;
  assign __muladd_madd_update_468 = _mul_21_stream_oready;

  madd_13
  __muladd_madd_468
  (
    .CLK(CLK),
    .update(__muladd_madd_update_468),
    .a(__delay_data_1869__delay_1868__delay_1867__variable_449),
    .b(__delay_data_1872__delay_1871__delay_1870__variable_450),
    .c(_cond_data_467),
    .d(__muladd_madd_odata_468)
  );

  reg [5-1:0] __delay_data_1876__delay_1875__delay_1874____variable_451;
  reg [5-1:0] __delay_data_1877__delay_1876__delay_1875____variable_451;
  reg [5-1:0] __delay_data_1878__delay_1877__delay_1876____variable_451;
  reg [5-1:0] __delay_data_1879__delay_1878__delay_1877____variable_451;
  reg signed [32-1:0] _sra_data_469;
  wire signed [32-1:0] mul_21_z_data;
  assign mul_21_z_data = _sra_data_469;
  wire signed [16-1:0] mul_22_x_data;
  wire signed [16-1:0] mul_22_y_data;
  wire [5-1:0] mul_22_rshift_data;
  reg __mul_22_stream_ivalid_1;
  reg __mul_22_stream_ivalid_2;
  reg __mul_22_stream_ivalid_3;
  reg __mul_22_stream_ivalid_4;
  reg __mul_22_stream_ivalid_5;
  reg __mul_22_stream_ivalid_6;
  reg __mul_22_stream_ivalid_7;
  reg __mul_22_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_473;
  reg [5-1:0] _minus_data_475;
  reg [1-1:0] _greatereq_data_486;
  reg signed [16-1:0] __delay_data_1886__variable_470;
  reg signed [16-1:0] __delay_data_1889__variable_471;
  reg [5-1:0] __delay_data_1892__variable_472;
  reg signed [34-1:0] _sll_data_477;
  reg [1-1:0] __delay_data_1883_greaterthan_473;
  reg [1-1:0] __delay_data_1884_greatereq_486;
  reg signed [16-1:0] __delay_data_1887__delay_1886__variable_470;
  reg signed [16-1:0] __delay_data_1890__delay_1889__variable_471;
  reg [5-1:0] __delay_data_1893__delay_1892__variable_472;
  reg signed [32-1:0] _cond_data_483;
  reg [1-1:0] __delay_data_1885__delay_1884_greatereq_486;
  reg signed [16-1:0] __delay_data_1888__delay_1887__delay_1886__variable_470;
  reg signed [16-1:0] __delay_data_1891__delay_1890__delay_1889__variable_471;
  reg [5-1:0] __delay_data_1894__delay_1893__delay_1892__variable_472;
  wire signed [16-1:0] _uminus_data_485;
  assign _uminus_data_485 = -_cond_data_483;
  wire signed [16-1:0] _cond_data_488;
  assign _cond_data_488 = (__delay_data_1885__delay_1884_greatereq_486)? _cond_data_483 : _uminus_data_485;
  wire signed [32-1:0] __muladd_madd_odata_489;
  reg signed [32-1:0] __muladd_madd_odata_reg_489;
  wire signed [32-1:0] __muladd_data_489;
  assign __muladd_data_489 = __muladd_madd_odata_reg_489;
  wire __muladd_madd_update_489;
  assign __muladd_madd_update_489 = _mul_22_stream_oready;

  madd_14
  __muladd_madd_489
  (
    .CLK(CLK),
    .update(__muladd_madd_update_489),
    .a(__delay_data_1888__delay_1887__delay_1886__variable_470),
    .b(__delay_data_1891__delay_1890__delay_1889__variable_471),
    .c(_cond_data_488),
    .d(__muladd_madd_odata_489)
  );

  reg [5-1:0] __delay_data_1895__delay_1894__delay_1893____variable_472;
  reg [5-1:0] __delay_data_1896__delay_1895__delay_1894____variable_472;
  reg [5-1:0] __delay_data_1897__delay_1896__delay_1895____variable_472;
  reg [5-1:0] __delay_data_1898__delay_1897__delay_1896____variable_472;
  reg signed [32-1:0] _sra_data_490;
  wire signed [32-1:0] mul_22_z_data;
  assign mul_22_z_data = _sra_data_490;
  wire signed [16-1:0] mul_23_x_data;
  wire signed [16-1:0] mul_23_y_data;
  wire [5-1:0] mul_23_rshift_data;
  reg __mul_23_stream_ivalid_1;
  reg __mul_23_stream_ivalid_2;
  reg __mul_23_stream_ivalid_3;
  reg __mul_23_stream_ivalid_4;
  reg __mul_23_stream_ivalid_5;
  reg __mul_23_stream_ivalid_6;
  reg __mul_23_stream_ivalid_7;
  reg __mul_23_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_494;
  reg [5-1:0] _minus_data_496;
  reg [1-1:0] _greatereq_data_507;
  reg signed [16-1:0] __delay_data_1905__variable_491;
  reg signed [16-1:0] __delay_data_1908__variable_492;
  reg [5-1:0] __delay_data_1911__variable_493;
  reg signed [34-1:0] _sll_data_498;
  reg [1-1:0] __delay_data_1902_greaterthan_494;
  reg [1-1:0] __delay_data_1903_greatereq_507;
  reg signed [16-1:0] __delay_data_1906__delay_1905__variable_491;
  reg signed [16-1:0] __delay_data_1909__delay_1908__variable_492;
  reg [5-1:0] __delay_data_1912__delay_1911__variable_493;
  reg signed [32-1:0] _cond_data_504;
  reg [1-1:0] __delay_data_1904__delay_1903_greatereq_507;
  reg signed [16-1:0] __delay_data_1907__delay_1906__delay_1905__variable_491;
  reg signed [16-1:0] __delay_data_1910__delay_1909__delay_1908__variable_492;
  reg [5-1:0] __delay_data_1913__delay_1912__delay_1911__variable_493;
  wire signed [16-1:0] _uminus_data_506;
  assign _uminus_data_506 = -_cond_data_504;
  wire signed [16-1:0] _cond_data_509;
  assign _cond_data_509 = (__delay_data_1904__delay_1903_greatereq_507)? _cond_data_504 : _uminus_data_506;
  wire signed [32-1:0] __muladd_madd_odata_510;
  reg signed [32-1:0] __muladd_madd_odata_reg_510;
  wire signed [32-1:0] __muladd_data_510;
  assign __muladd_data_510 = __muladd_madd_odata_reg_510;
  wire __muladd_madd_update_510;
  assign __muladd_madd_update_510 = _mul_23_stream_oready;

  madd_15
  __muladd_madd_510
  (
    .CLK(CLK),
    .update(__muladd_madd_update_510),
    .a(__delay_data_1907__delay_1906__delay_1905__variable_491),
    .b(__delay_data_1910__delay_1909__delay_1908__variable_492),
    .c(_cond_data_509),
    .d(__muladd_madd_odata_510)
  );

  reg [5-1:0] __delay_data_1914__delay_1913__delay_1912____variable_493;
  reg [5-1:0] __delay_data_1915__delay_1914__delay_1913____variable_493;
  reg [5-1:0] __delay_data_1916__delay_1915__delay_1914____variable_493;
  reg [5-1:0] __delay_data_1917__delay_1916__delay_1915____variable_493;
  reg signed [32-1:0] _sra_data_511;
  wire signed [32-1:0] mul_23_z_data;
  assign mul_23_z_data = _sra_data_511;
  wire signed [16-1:0] mul_24_x_data;
  wire signed [16-1:0] mul_24_y_data;
  wire [5-1:0] mul_24_rshift_data;
  reg __mul_24_stream_ivalid_1;
  reg __mul_24_stream_ivalid_2;
  reg __mul_24_stream_ivalid_3;
  reg __mul_24_stream_ivalid_4;
  reg __mul_24_stream_ivalid_5;
  reg __mul_24_stream_ivalid_6;
  reg __mul_24_stream_ivalid_7;
  reg __mul_24_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_515;
  reg [5-1:0] _minus_data_517;
  reg [1-1:0] _greatereq_data_528;
  reg signed [16-1:0] __delay_data_1924__variable_512;
  reg signed [16-1:0] __delay_data_1927__variable_513;
  reg [5-1:0] __delay_data_1930__variable_514;
  reg signed [34-1:0] _sll_data_519;
  reg [1-1:0] __delay_data_1921_greaterthan_515;
  reg [1-1:0] __delay_data_1922_greatereq_528;
  reg signed [16-1:0] __delay_data_1925__delay_1924__variable_512;
  reg signed [16-1:0] __delay_data_1928__delay_1927__variable_513;
  reg [5-1:0] __delay_data_1931__delay_1930__variable_514;
  reg signed [32-1:0] _cond_data_525;
  reg [1-1:0] __delay_data_1923__delay_1922_greatereq_528;
  reg signed [16-1:0] __delay_data_1926__delay_1925__delay_1924__variable_512;
  reg signed [16-1:0] __delay_data_1929__delay_1928__delay_1927__variable_513;
  reg [5-1:0] __delay_data_1932__delay_1931__delay_1930__variable_514;
  wire signed [16-1:0] _uminus_data_527;
  assign _uminus_data_527 = -_cond_data_525;
  wire signed [16-1:0] _cond_data_530;
  assign _cond_data_530 = (__delay_data_1923__delay_1922_greatereq_528)? _cond_data_525 : _uminus_data_527;
  wire signed [32-1:0] __muladd_madd_odata_531;
  reg signed [32-1:0] __muladd_madd_odata_reg_531;
  wire signed [32-1:0] __muladd_data_531;
  assign __muladd_data_531 = __muladd_madd_odata_reg_531;
  wire __muladd_madd_update_531;
  assign __muladd_madd_update_531 = _mul_24_stream_oready;

  madd_16
  __muladd_madd_531
  (
    .CLK(CLK),
    .update(__muladd_madd_update_531),
    .a(__delay_data_1926__delay_1925__delay_1924__variable_512),
    .b(__delay_data_1929__delay_1928__delay_1927__variable_513),
    .c(_cond_data_530),
    .d(__muladd_madd_odata_531)
  );

  reg [5-1:0] __delay_data_1933__delay_1932__delay_1931____variable_514;
  reg [5-1:0] __delay_data_1934__delay_1933__delay_1932____variable_514;
  reg [5-1:0] __delay_data_1935__delay_1934__delay_1933____variable_514;
  reg [5-1:0] __delay_data_1936__delay_1935__delay_1934____variable_514;
  reg signed [32-1:0] _sra_data_532;
  wire signed [32-1:0] mul_24_z_data;
  assign mul_24_z_data = _sra_data_532;
  wire signed [16-1:0] mul_25_x_data;
  wire signed [16-1:0] mul_25_y_data;
  wire [5-1:0] mul_25_rshift_data;
  reg __mul_25_stream_ivalid_1;
  reg __mul_25_stream_ivalid_2;
  reg __mul_25_stream_ivalid_3;
  reg __mul_25_stream_ivalid_4;
  reg __mul_25_stream_ivalid_5;
  reg __mul_25_stream_ivalid_6;
  reg __mul_25_stream_ivalid_7;
  reg __mul_25_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_536;
  reg [5-1:0] _minus_data_538;
  reg [1-1:0] _greatereq_data_549;
  reg signed [16-1:0] __delay_data_1943__variable_533;
  reg signed [16-1:0] __delay_data_1946__variable_534;
  reg [5-1:0] __delay_data_1949__variable_535;
  reg signed [34-1:0] _sll_data_540;
  reg [1-1:0] __delay_data_1940_greaterthan_536;
  reg [1-1:0] __delay_data_1941_greatereq_549;
  reg signed [16-1:0] __delay_data_1944__delay_1943__variable_533;
  reg signed [16-1:0] __delay_data_1947__delay_1946__variable_534;
  reg [5-1:0] __delay_data_1950__delay_1949__variable_535;
  reg signed [32-1:0] _cond_data_546;
  reg [1-1:0] __delay_data_1942__delay_1941_greatereq_549;
  reg signed [16-1:0] __delay_data_1945__delay_1944__delay_1943__variable_533;
  reg signed [16-1:0] __delay_data_1948__delay_1947__delay_1946__variable_534;
  reg [5-1:0] __delay_data_1951__delay_1950__delay_1949__variable_535;
  wire signed [16-1:0] _uminus_data_548;
  assign _uminus_data_548 = -_cond_data_546;
  wire signed [16-1:0] _cond_data_551;
  assign _cond_data_551 = (__delay_data_1942__delay_1941_greatereq_549)? _cond_data_546 : _uminus_data_548;
  wire signed [32-1:0] __muladd_madd_odata_552;
  reg signed [32-1:0] __muladd_madd_odata_reg_552;
  wire signed [32-1:0] __muladd_data_552;
  assign __muladd_data_552 = __muladd_madd_odata_reg_552;
  wire __muladd_madd_update_552;
  assign __muladd_madd_update_552 = _mul_25_stream_oready;

  madd_17
  __muladd_madd_552
  (
    .CLK(CLK),
    .update(__muladd_madd_update_552),
    .a(__delay_data_1945__delay_1944__delay_1943__variable_533),
    .b(__delay_data_1948__delay_1947__delay_1946__variable_534),
    .c(_cond_data_551),
    .d(__muladd_madd_odata_552)
  );

  reg [5-1:0] __delay_data_1952__delay_1951__delay_1950____variable_535;
  reg [5-1:0] __delay_data_1953__delay_1952__delay_1951____variable_535;
  reg [5-1:0] __delay_data_1954__delay_1953__delay_1952____variable_535;
  reg [5-1:0] __delay_data_1955__delay_1954__delay_1953____variable_535;
  reg signed [32-1:0] _sra_data_553;
  wire signed [32-1:0] mul_25_z_data;
  assign mul_25_z_data = _sra_data_553;
  wire signed [64-1:0] add_tree_4_var0_data;
  wire signed [64-1:0] add_tree_4_var1_data;
  wire signed [64-1:0] add_tree_4_var2_data;
  wire signed [64-1:0] add_tree_4_var3_data;
  wire signed [64-1:0] add_tree_4_var4_data;
  wire signed [64-1:0] add_tree_4_var5_data;
  wire signed [64-1:0] add_tree_4_var6_data;
  wire signed [64-1:0] add_tree_4_var7_data;
  wire signed [64-1:0] add_tree_4_var8_data;
  wire signed [64-1:0] add_tree_4_var9_data;
  wire signed [64-1:0] add_tree_4_var10_data;
  wire signed [64-1:0] add_tree_4_var11_data;
  wire signed [64-1:0] add_tree_4_var12_data;
  wire signed [64-1:0] add_tree_4_var13_data;
  wire signed [64-1:0] add_tree_4_var14_data;
  wire signed [64-1:0] add_tree_4_var15_data;
  wire signed [64-1:0] add_tree_4_var16_data;
  wire signed [64-1:0] add_tree_4_var17_data;
  reg __add_tree_4_stream_ivalid_1;
  reg __add_tree_4_stream_ivalid_2;
  reg __add_tree_4_stream_ivalid_3;
  reg signed [64-1:0] __plusn_data_71;
  reg signed [64-1:0] __plusn_data_72;
  reg signed [64-1:0] __plusn_data_73;
  reg signed [64-1:0] __plusn_data_75;
  reg signed [64-1:0] __plusn_data_76;
  reg signed [64-1:0] __plusn_data_77;
  reg signed [64-1:0] __plusn_data_74;
  reg signed [64-1:0] __plusn_data_78;
  reg signed [64-1:0] __plusn_data_79;
  wire signed [64-1:0] add_tree_4_sum_data;
  assign add_tree_4_sum_data = __plusn_data_79;
  wire signed [64-1:0] acc_0_x_data;
  wire [7-1:0] acc_0_rshift_data;
  wire [32-1:0] acc_0_size_data;
  wire [1-1:0] acc_0__reduce_reset_data;
  reg __acc_0_stream_ivalid_1;
  reg __acc_0_stream_ivalid_2;
  reg __acc_0_stream_ivalid_3;
  reg __acc_0_stream_ivalid_4;
  reg __acc_0_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_3;
  reg [7-1:0] _minus_data_5;
  reg signed [64-1:0] _reduceadd_data_16;
  reg [33-1:0] _reduceadd_count_16;
  reg _reduceadd_prev_count_max_16;
  wire _reduceadd_reset_cond_16;
  assign _reduceadd_reset_cond_16 = acc_0__reduce_reset_data || _reduceadd_prev_count_max_16;
  wire [33-1:0] _reduceadd_current_count_16;
  assign _reduceadd_current_count_16 = (_reduceadd_reset_cond_16)? 0 : _reduceadd_count_16;
  wire signed [64-1:0] _reduceadd_current_data_16;
  assign _reduceadd_current_data_16 = (_reduceadd_reset_cond_16)? 1'sd0 : _reduceadd_data_16;
  reg [1-1:0] _pulse_data_18;
  reg [33-1:0] _pulse_count_18;
  reg _pulse_prev_count_max_18;
  wire _pulse_reset_cond_18;
  assign _pulse_reset_cond_18 = acc_0__reduce_reset_data || _pulse_prev_count_max_18;
  wire [33-1:0] _pulse_current_count_18;
  assign _pulse_current_count_18 = (_pulse_reset_cond_18)? 0 : _pulse_count_18;
  wire [1-1:0] _pulse_current_data_18;
  assign _pulse_current_data_18 = (_pulse_reset_cond_18)? 1'sd0 : _pulse_data_18;
  reg [7-1:0] __delay_data_1964__variable_1;
  reg signed [130-1:0] _sll_data_7;
  reg [1-1:0] __delay_data_1961_greaterthan_3;
  reg signed [64-1:0] __delay_data_1962_reduceadd_16;
  reg [7-1:0] __delay_data_1965__delay_1964__variable_1;
  reg [1-1:0] __delay_data_1968_pulse_18;
  reg signed [64-1:0] _cond_data_13;
  reg signed [64-1:0] __delay_data_1963__delay_1962_reduceadd_16;
  reg [7-1:0] __delay_data_1966__delay_1965__delay_1964__variable_1;
  reg [1-1:0] __delay_data_1969__delay_1968_pulse_18;
  reg signed [64-1:0] _plus_data_20;
  reg [7-1:0] __delay_data_1967__delay_1966__delay_1965____variable_1;
  reg [1-1:0] __delay_data_1970__delay_1969__delay_1968_pulse_18;
  reg signed [64-1:0] _sra_data_21;
  reg [1-1:0] __delay_data_1971__delay_1970__delay_1969__delay_1968_pulse_18;
  wire signed [64-1:0] acc_0_sum_data;
  assign acc_0_sum_data = _sra_data_21;
  wire [1-1:0] acc_0_valid_data;
  assign acc_0_valid_data = __delay_data_1971__delay_1970__delay_1969__delay_1968_pulse_18;
  wire signed [64-1:0] mul_rshift_round_clip_6_x_data;
  wire signed [16-1:0] mul_rshift_round_clip_6_y_data;
  wire [7-1:0] mul_rshift_round_clip_6_rshift_data;
  reg __mul_rshift_round_clip_6_stream_ivalid_1;
  reg __mul_rshift_round_clip_6_stream_ivalid_2;
  reg __mul_rshift_round_clip_6_stream_ivalid_3;
  reg __mul_rshift_round_clip_6_stream_ivalid_4;
  reg __mul_rshift_round_clip_6_stream_ivalid_5;
  reg __mul_rshift_round_clip_6_stream_ivalid_6;
  reg __mul_rshift_round_clip_6_stream_ivalid_7;
  reg __mul_rshift_round_clip_6_stream_ivalid_8;
  wire signed [80-1:0] _times_mul_odata_111;
  reg signed [80-1:0] _times_mul_odata_reg_111;
  wire signed [80-1:0] _times_data_111;
  assign _times_data_111 = _times_mul_odata_reg_111;
  wire _times_mul_update_111;
  assign _times_mul_update_111 = _mul_rshift_round_clip_6_stream_oready;

  multiplier_0
  _times_mul_111
  (
    .CLK(CLK),
    .update(_times_mul_update_111),
    .a(mul_rshift_round_clip_6_x_data),
    .b(mul_rshift_round_clip_6_y_data),
    .c(_times_mul_odata_111)
  );

  wire [7-1:0] _minus_data_114;
  assign _minus_data_114 = mul_rshift_round_clip_6_rshift_data - 2'sd1;
  wire signed [130-1:0] _sll_data_117;
  assign _sll_data_117 = 2'sd1 << _minus_data_114;
  wire [1-1:0] _eq_data_129;
  assign _eq_data_129 = mul_rshift_round_clip_6_rshift_data == 1'sd0;
  reg signed [130-1:0] __delay_data_1977_sll_117;
  reg [7-1:0] __delay_data_1981__variable_110;
  reg [1-1:0] __delay_data_1985_eq_129;
  reg signed [130-1:0] __delay_data_1978__delay_1977_sll_117;
  reg [7-1:0] __delay_data_1982__delay_1981__variable_110;
  reg [1-1:0] __delay_data_1986__delay_1985_eq_129;
  reg signed [130-1:0] __delay_data_1979__delay_1978__delay_1977_sll_117;
  reg [7-1:0] __delay_data_1983__delay_1982__delay_1981__variable_110;
  reg [1-1:0] __delay_data_1987__delay_1986__delay_1985_eq_129;
  reg signed [130-1:0] __delay_data_1980__delay_1979__delay_1978__delay_1977_sll_117;
  reg [7-1:0] __delay_data_1984__delay_1983__delay_1982____variable_110;
  reg [1-1:0] __delay_data_1988__delay_1987__delay_1986__delay_1985_eq_129;
  wire [1-1:0] _pointer_data_112;
  assign _pointer_data_112 = _times_data_111[8'sd79];
  wire signed [2-1:0] _cond_data_124;
  assign _cond_data_124 = (_pointer_data_112)? -2'sd1 : 1'sd0;
  wire signed [81-1:0] _plus_data_125;
  assign _plus_data_125 = _times_data_111 + __delay_data_1980__delay_1979__delay_1978__delay_1977_sll_117;
  wire signed [81-1:0] _plus_data_126;
  assign _plus_data_126 = _plus_data_125 + _cond_data_124;
  wire signed [80-1:0] _sra_data_127;
  assign _sra_data_127 = _plus_data_126 >>> __delay_data_1984__delay_1983__delay_1982____variable_110;
  reg signed [80-1:0] _cond_data_130;
  reg [1-1:0] _greaterthan_data_131;
  reg [1-1:0] _lessthan_data_135;
  reg [1-1:0] _greatereq_data_139;
  reg signed [80-1:0] __delay_data_1989_cond_130;
  reg signed [80-1:0] _cond_data_133;
  reg signed [80-1:0] _cond_data_137;
  reg [1-1:0] __delay_data_1990_greatereq_139;
  reg signed [16-1:0] _cond_data_141;
  wire signed [16-1:0] mul_rshift_round_clip_6_z_data;
  assign mul_rshift_round_clip_6_z_data = _cond_data_141;
  wire signed [16-1:0] mul_26_x_data;
  wire signed [16-1:0] mul_26_y_data;
  wire [5-1:0] mul_26_rshift_data;
  reg __mul_26_stream_ivalid_1;
  reg __mul_26_stream_ivalid_2;
  reg __mul_26_stream_ivalid_3;
  reg __mul_26_stream_ivalid_4;
  reg __mul_26_stream_ivalid_5;
  reg __mul_26_stream_ivalid_6;
  reg __mul_26_stream_ivalid_7;
  reg __mul_26_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_557;
  reg [5-1:0] _minus_data_559;
  reg [1-1:0] _greatereq_data_570;
  reg signed [16-1:0] __delay_data_2020__variable_554;
  reg signed [16-1:0] __delay_data_2023__variable_555;
  reg [5-1:0] __delay_data_2026__variable_556;
  reg signed [34-1:0] _sll_data_561;
  reg [1-1:0] __delay_data_2017_greaterthan_557;
  reg [1-1:0] __delay_data_2018_greatereq_570;
  reg signed [16-1:0] __delay_data_2021__delay_2020__variable_554;
  reg signed [16-1:0] __delay_data_2024__delay_2023__variable_555;
  reg [5-1:0] __delay_data_2027__delay_2026__variable_556;
  reg signed [32-1:0] _cond_data_567;
  reg [1-1:0] __delay_data_2019__delay_2018_greatereq_570;
  reg signed [16-1:0] __delay_data_2022__delay_2021__delay_2020__variable_554;
  reg signed [16-1:0] __delay_data_2025__delay_2024__delay_2023__variable_555;
  reg [5-1:0] __delay_data_2028__delay_2027__delay_2026__variable_556;
  wire signed [16-1:0] _uminus_data_569;
  assign _uminus_data_569 = -_cond_data_567;
  wire signed [16-1:0] _cond_data_572;
  assign _cond_data_572 = (__delay_data_2019__delay_2018_greatereq_570)? _cond_data_567 : _uminus_data_569;
  wire signed [32-1:0] __muladd_madd_odata_573;
  reg signed [32-1:0] __muladd_madd_odata_reg_573;
  wire signed [32-1:0] __muladd_data_573;
  assign __muladd_data_573 = __muladd_madd_odata_reg_573;
  wire __muladd_madd_update_573;
  assign __muladd_madd_update_573 = _mul_26_stream_oready;

  madd_18
  __muladd_madd_573
  (
    .CLK(CLK),
    .update(__muladd_madd_update_573),
    .a(__delay_data_2022__delay_2021__delay_2020__variable_554),
    .b(__delay_data_2025__delay_2024__delay_2023__variable_555),
    .c(_cond_data_572),
    .d(__muladd_madd_odata_573)
  );

  reg [5-1:0] __delay_data_2029__delay_2028__delay_2027____variable_556;
  reg [5-1:0] __delay_data_2030__delay_2029__delay_2028____variable_556;
  reg [5-1:0] __delay_data_2031__delay_2030__delay_2029____variable_556;
  reg [5-1:0] __delay_data_2032__delay_2031__delay_2030____variable_556;
  reg signed [32-1:0] _sra_data_574;
  wire signed [32-1:0] mul_26_z_data;
  assign mul_26_z_data = _sra_data_574;
  wire signed [16-1:0] mul_27_x_data;
  wire signed [16-1:0] mul_27_y_data;
  wire [5-1:0] mul_27_rshift_data;
  reg __mul_27_stream_ivalid_1;
  reg __mul_27_stream_ivalid_2;
  reg __mul_27_stream_ivalid_3;
  reg __mul_27_stream_ivalid_4;
  reg __mul_27_stream_ivalid_5;
  reg __mul_27_stream_ivalid_6;
  reg __mul_27_stream_ivalid_7;
  reg __mul_27_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_578;
  reg [5-1:0] _minus_data_580;
  reg [1-1:0] _greatereq_data_591;
  reg signed [16-1:0] __delay_data_2039__variable_575;
  reg signed [16-1:0] __delay_data_2042__variable_576;
  reg [5-1:0] __delay_data_2045__variable_577;
  reg signed [34-1:0] _sll_data_582;
  reg [1-1:0] __delay_data_2036_greaterthan_578;
  reg [1-1:0] __delay_data_2037_greatereq_591;
  reg signed [16-1:0] __delay_data_2040__delay_2039__variable_575;
  reg signed [16-1:0] __delay_data_2043__delay_2042__variable_576;
  reg [5-1:0] __delay_data_2046__delay_2045__variable_577;
  reg signed [32-1:0] _cond_data_588;
  reg [1-1:0] __delay_data_2038__delay_2037_greatereq_591;
  reg signed [16-1:0] __delay_data_2041__delay_2040__delay_2039__variable_575;
  reg signed [16-1:0] __delay_data_2044__delay_2043__delay_2042__variable_576;
  reg [5-1:0] __delay_data_2047__delay_2046__delay_2045__variable_577;
  wire signed [16-1:0] _uminus_data_590;
  assign _uminus_data_590 = -_cond_data_588;
  wire signed [16-1:0] _cond_data_593;
  assign _cond_data_593 = (__delay_data_2038__delay_2037_greatereq_591)? _cond_data_588 : _uminus_data_590;
  wire signed [32-1:0] __muladd_madd_odata_594;
  reg signed [32-1:0] __muladd_madd_odata_reg_594;
  wire signed [32-1:0] __muladd_data_594;
  assign __muladd_data_594 = __muladd_madd_odata_reg_594;
  wire __muladd_madd_update_594;
  assign __muladd_madd_update_594 = _mul_27_stream_oready;

  madd_19
  __muladd_madd_594
  (
    .CLK(CLK),
    .update(__muladd_madd_update_594),
    .a(__delay_data_2041__delay_2040__delay_2039__variable_575),
    .b(__delay_data_2044__delay_2043__delay_2042__variable_576),
    .c(_cond_data_593),
    .d(__muladd_madd_odata_594)
  );

  reg [5-1:0] __delay_data_2048__delay_2047__delay_2046____variable_577;
  reg [5-1:0] __delay_data_2049__delay_2048__delay_2047____variable_577;
  reg [5-1:0] __delay_data_2050__delay_2049__delay_2048____variable_577;
  reg [5-1:0] __delay_data_2051__delay_2050__delay_2049____variable_577;
  reg signed [32-1:0] _sra_data_595;
  wire signed [32-1:0] mul_27_z_data;
  assign mul_27_z_data = _sra_data_595;
  wire signed [16-1:0] mul_28_x_data;
  wire signed [16-1:0] mul_28_y_data;
  wire [5-1:0] mul_28_rshift_data;
  reg __mul_28_stream_ivalid_1;
  reg __mul_28_stream_ivalid_2;
  reg __mul_28_stream_ivalid_3;
  reg __mul_28_stream_ivalid_4;
  reg __mul_28_stream_ivalid_5;
  reg __mul_28_stream_ivalid_6;
  reg __mul_28_stream_ivalid_7;
  reg __mul_28_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_599;
  reg [5-1:0] _minus_data_601;
  reg [1-1:0] _greatereq_data_612;
  reg signed [16-1:0] __delay_data_2058__variable_596;
  reg signed [16-1:0] __delay_data_2061__variable_597;
  reg [5-1:0] __delay_data_2064__variable_598;
  reg signed [34-1:0] _sll_data_603;
  reg [1-1:0] __delay_data_2055_greaterthan_599;
  reg [1-1:0] __delay_data_2056_greatereq_612;
  reg signed [16-1:0] __delay_data_2059__delay_2058__variable_596;
  reg signed [16-1:0] __delay_data_2062__delay_2061__variable_597;
  reg [5-1:0] __delay_data_2065__delay_2064__variable_598;
  reg signed [32-1:0] _cond_data_609;
  reg [1-1:0] __delay_data_2057__delay_2056_greatereq_612;
  reg signed [16-1:0] __delay_data_2060__delay_2059__delay_2058__variable_596;
  reg signed [16-1:0] __delay_data_2063__delay_2062__delay_2061__variable_597;
  reg [5-1:0] __delay_data_2066__delay_2065__delay_2064__variable_598;
  wire signed [16-1:0] _uminus_data_611;
  assign _uminus_data_611 = -_cond_data_609;
  wire signed [16-1:0] _cond_data_614;
  assign _cond_data_614 = (__delay_data_2057__delay_2056_greatereq_612)? _cond_data_609 : _uminus_data_611;
  wire signed [32-1:0] __muladd_madd_odata_615;
  reg signed [32-1:0] __muladd_madd_odata_reg_615;
  wire signed [32-1:0] __muladd_data_615;
  assign __muladd_data_615 = __muladd_madd_odata_reg_615;
  wire __muladd_madd_update_615;
  assign __muladd_madd_update_615 = _mul_28_stream_oready;

  madd_20
  __muladd_madd_615
  (
    .CLK(CLK),
    .update(__muladd_madd_update_615),
    .a(__delay_data_2060__delay_2059__delay_2058__variable_596),
    .b(__delay_data_2063__delay_2062__delay_2061__variable_597),
    .c(_cond_data_614),
    .d(__muladd_madd_odata_615)
  );

  reg [5-1:0] __delay_data_2067__delay_2066__delay_2065____variable_598;
  reg [5-1:0] __delay_data_2068__delay_2067__delay_2066____variable_598;
  reg [5-1:0] __delay_data_2069__delay_2068__delay_2067____variable_598;
  reg [5-1:0] __delay_data_2070__delay_2069__delay_2068____variable_598;
  reg signed [32-1:0] _sra_data_616;
  wire signed [32-1:0] mul_28_z_data;
  assign mul_28_z_data = _sra_data_616;
  wire signed [16-1:0] mul_29_x_data;
  wire signed [16-1:0] mul_29_y_data;
  wire [5-1:0] mul_29_rshift_data;
  reg __mul_29_stream_ivalid_1;
  reg __mul_29_stream_ivalid_2;
  reg __mul_29_stream_ivalid_3;
  reg __mul_29_stream_ivalid_4;
  reg __mul_29_stream_ivalid_5;
  reg __mul_29_stream_ivalid_6;
  reg __mul_29_stream_ivalid_7;
  reg __mul_29_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_620;
  reg [5-1:0] _minus_data_622;
  reg [1-1:0] _greatereq_data_633;
  reg signed [16-1:0] __delay_data_2077__variable_617;
  reg signed [16-1:0] __delay_data_2080__variable_618;
  reg [5-1:0] __delay_data_2083__variable_619;
  reg signed [34-1:0] _sll_data_624;
  reg [1-1:0] __delay_data_2074_greaterthan_620;
  reg [1-1:0] __delay_data_2075_greatereq_633;
  reg signed [16-1:0] __delay_data_2078__delay_2077__variable_617;
  reg signed [16-1:0] __delay_data_2081__delay_2080__variable_618;
  reg [5-1:0] __delay_data_2084__delay_2083__variable_619;
  reg signed [32-1:0] _cond_data_630;
  reg [1-1:0] __delay_data_2076__delay_2075_greatereq_633;
  reg signed [16-1:0] __delay_data_2079__delay_2078__delay_2077__variable_617;
  reg signed [16-1:0] __delay_data_2082__delay_2081__delay_2080__variable_618;
  reg [5-1:0] __delay_data_2085__delay_2084__delay_2083__variable_619;
  wire signed [16-1:0] _uminus_data_632;
  assign _uminus_data_632 = -_cond_data_630;
  wire signed [16-1:0] _cond_data_635;
  assign _cond_data_635 = (__delay_data_2076__delay_2075_greatereq_633)? _cond_data_630 : _uminus_data_632;
  wire signed [32-1:0] __muladd_madd_odata_636;
  reg signed [32-1:0] __muladd_madd_odata_reg_636;
  wire signed [32-1:0] __muladd_data_636;
  assign __muladd_data_636 = __muladd_madd_odata_reg_636;
  wire __muladd_madd_update_636;
  assign __muladd_madd_update_636 = _mul_29_stream_oready;

  madd_21
  __muladd_madd_636
  (
    .CLK(CLK),
    .update(__muladd_madd_update_636),
    .a(__delay_data_2079__delay_2078__delay_2077__variable_617),
    .b(__delay_data_2082__delay_2081__delay_2080__variable_618),
    .c(_cond_data_635),
    .d(__muladd_madd_odata_636)
  );

  reg [5-1:0] __delay_data_2086__delay_2085__delay_2084____variable_619;
  reg [5-1:0] __delay_data_2087__delay_2086__delay_2085____variable_619;
  reg [5-1:0] __delay_data_2088__delay_2087__delay_2086____variable_619;
  reg [5-1:0] __delay_data_2089__delay_2088__delay_2087____variable_619;
  reg signed [32-1:0] _sra_data_637;
  wire signed [32-1:0] mul_29_z_data;
  assign mul_29_z_data = _sra_data_637;
  wire signed [16-1:0] mul_30_x_data;
  wire signed [16-1:0] mul_30_y_data;
  wire [5-1:0] mul_30_rshift_data;
  reg __mul_30_stream_ivalid_1;
  reg __mul_30_stream_ivalid_2;
  reg __mul_30_stream_ivalid_3;
  reg __mul_30_stream_ivalid_4;
  reg __mul_30_stream_ivalid_5;
  reg __mul_30_stream_ivalid_6;
  reg __mul_30_stream_ivalid_7;
  reg __mul_30_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_641;
  reg [5-1:0] _minus_data_643;
  reg [1-1:0] _greatereq_data_654;
  reg signed [16-1:0] __delay_data_2096__variable_638;
  reg signed [16-1:0] __delay_data_2099__variable_639;
  reg [5-1:0] __delay_data_2102__variable_640;
  reg signed [34-1:0] _sll_data_645;
  reg [1-1:0] __delay_data_2093_greaterthan_641;
  reg [1-1:0] __delay_data_2094_greatereq_654;
  reg signed [16-1:0] __delay_data_2097__delay_2096__variable_638;
  reg signed [16-1:0] __delay_data_2100__delay_2099__variable_639;
  reg [5-1:0] __delay_data_2103__delay_2102__variable_640;
  reg signed [32-1:0] _cond_data_651;
  reg [1-1:0] __delay_data_2095__delay_2094_greatereq_654;
  reg signed [16-1:0] __delay_data_2098__delay_2097__delay_2096__variable_638;
  reg signed [16-1:0] __delay_data_2101__delay_2100__delay_2099__variable_639;
  reg [5-1:0] __delay_data_2104__delay_2103__delay_2102__variable_640;
  wire signed [16-1:0] _uminus_data_653;
  assign _uminus_data_653 = -_cond_data_651;
  wire signed [16-1:0] _cond_data_656;
  assign _cond_data_656 = (__delay_data_2095__delay_2094_greatereq_654)? _cond_data_651 : _uminus_data_653;
  wire signed [32-1:0] __muladd_madd_odata_657;
  reg signed [32-1:0] __muladd_madd_odata_reg_657;
  wire signed [32-1:0] __muladd_data_657;
  assign __muladd_data_657 = __muladd_madd_odata_reg_657;
  wire __muladd_madd_update_657;
  assign __muladd_madd_update_657 = _mul_30_stream_oready;

  madd_22
  __muladd_madd_657
  (
    .CLK(CLK),
    .update(__muladd_madd_update_657),
    .a(__delay_data_2098__delay_2097__delay_2096__variable_638),
    .b(__delay_data_2101__delay_2100__delay_2099__variable_639),
    .c(_cond_data_656),
    .d(__muladd_madd_odata_657)
  );

  reg [5-1:0] __delay_data_2105__delay_2104__delay_2103____variable_640;
  reg [5-1:0] __delay_data_2106__delay_2105__delay_2104____variable_640;
  reg [5-1:0] __delay_data_2107__delay_2106__delay_2105____variable_640;
  reg [5-1:0] __delay_data_2108__delay_2107__delay_2106____variable_640;
  reg signed [32-1:0] _sra_data_658;
  wire signed [32-1:0] mul_30_z_data;
  assign mul_30_z_data = _sra_data_658;
  wire signed [16-1:0] mul_31_x_data;
  wire signed [16-1:0] mul_31_y_data;
  wire [5-1:0] mul_31_rshift_data;
  reg __mul_31_stream_ivalid_1;
  reg __mul_31_stream_ivalid_2;
  reg __mul_31_stream_ivalid_3;
  reg __mul_31_stream_ivalid_4;
  reg __mul_31_stream_ivalid_5;
  reg __mul_31_stream_ivalid_6;
  reg __mul_31_stream_ivalid_7;
  reg __mul_31_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_662;
  reg [5-1:0] _minus_data_664;
  reg [1-1:0] _greatereq_data_675;
  reg signed [16-1:0] __delay_data_2115__variable_659;
  reg signed [16-1:0] __delay_data_2118__variable_660;
  reg [5-1:0] __delay_data_2121__variable_661;
  reg signed [34-1:0] _sll_data_666;
  reg [1-1:0] __delay_data_2112_greaterthan_662;
  reg [1-1:0] __delay_data_2113_greatereq_675;
  reg signed [16-1:0] __delay_data_2116__delay_2115__variable_659;
  reg signed [16-1:0] __delay_data_2119__delay_2118__variable_660;
  reg [5-1:0] __delay_data_2122__delay_2121__variable_661;
  reg signed [32-1:0] _cond_data_672;
  reg [1-1:0] __delay_data_2114__delay_2113_greatereq_675;
  reg signed [16-1:0] __delay_data_2117__delay_2116__delay_2115__variable_659;
  reg signed [16-1:0] __delay_data_2120__delay_2119__delay_2118__variable_660;
  reg [5-1:0] __delay_data_2123__delay_2122__delay_2121__variable_661;
  wire signed [16-1:0] _uminus_data_674;
  assign _uminus_data_674 = -_cond_data_672;
  wire signed [16-1:0] _cond_data_677;
  assign _cond_data_677 = (__delay_data_2114__delay_2113_greatereq_675)? _cond_data_672 : _uminus_data_674;
  wire signed [32-1:0] __muladd_madd_odata_678;
  reg signed [32-1:0] __muladd_madd_odata_reg_678;
  wire signed [32-1:0] __muladd_data_678;
  assign __muladd_data_678 = __muladd_madd_odata_reg_678;
  wire __muladd_madd_update_678;
  assign __muladd_madd_update_678 = _mul_31_stream_oready;

  madd_23
  __muladd_madd_678
  (
    .CLK(CLK),
    .update(__muladd_madd_update_678),
    .a(__delay_data_2117__delay_2116__delay_2115__variable_659),
    .b(__delay_data_2120__delay_2119__delay_2118__variable_660),
    .c(_cond_data_677),
    .d(__muladd_madd_odata_678)
  );

  reg [5-1:0] __delay_data_2124__delay_2123__delay_2122____variable_661;
  reg [5-1:0] __delay_data_2125__delay_2124__delay_2123____variable_661;
  reg [5-1:0] __delay_data_2126__delay_2125__delay_2124____variable_661;
  reg [5-1:0] __delay_data_2127__delay_2126__delay_2125____variable_661;
  reg signed [32-1:0] _sra_data_679;
  wire signed [32-1:0] mul_31_z_data;
  assign mul_31_z_data = _sra_data_679;
  wire signed [16-1:0] mul_32_x_data;
  wire signed [16-1:0] mul_32_y_data;
  wire [5-1:0] mul_32_rshift_data;
  reg __mul_32_stream_ivalid_1;
  reg __mul_32_stream_ivalid_2;
  reg __mul_32_stream_ivalid_3;
  reg __mul_32_stream_ivalid_4;
  reg __mul_32_stream_ivalid_5;
  reg __mul_32_stream_ivalid_6;
  reg __mul_32_stream_ivalid_7;
  reg __mul_32_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_683;
  reg [5-1:0] _minus_data_685;
  reg [1-1:0] _greatereq_data_696;
  reg signed [16-1:0] __delay_data_2134__variable_680;
  reg signed [16-1:0] __delay_data_2137__variable_681;
  reg [5-1:0] __delay_data_2140__variable_682;
  reg signed [34-1:0] _sll_data_687;
  reg [1-1:0] __delay_data_2131_greaterthan_683;
  reg [1-1:0] __delay_data_2132_greatereq_696;
  reg signed [16-1:0] __delay_data_2135__delay_2134__variable_680;
  reg signed [16-1:0] __delay_data_2138__delay_2137__variable_681;
  reg [5-1:0] __delay_data_2141__delay_2140__variable_682;
  reg signed [32-1:0] _cond_data_693;
  reg [1-1:0] __delay_data_2133__delay_2132_greatereq_696;
  reg signed [16-1:0] __delay_data_2136__delay_2135__delay_2134__variable_680;
  reg signed [16-1:0] __delay_data_2139__delay_2138__delay_2137__variable_681;
  reg [5-1:0] __delay_data_2142__delay_2141__delay_2140__variable_682;
  wire signed [16-1:0] _uminus_data_695;
  assign _uminus_data_695 = -_cond_data_693;
  wire signed [16-1:0] _cond_data_698;
  assign _cond_data_698 = (__delay_data_2133__delay_2132_greatereq_696)? _cond_data_693 : _uminus_data_695;
  wire signed [32-1:0] __muladd_madd_odata_699;
  reg signed [32-1:0] __muladd_madd_odata_reg_699;
  wire signed [32-1:0] __muladd_data_699;
  assign __muladd_data_699 = __muladd_madd_odata_reg_699;
  wire __muladd_madd_update_699;
  assign __muladd_madd_update_699 = _mul_32_stream_oready;

  madd_24
  __muladd_madd_699
  (
    .CLK(CLK),
    .update(__muladd_madd_update_699),
    .a(__delay_data_2136__delay_2135__delay_2134__variable_680),
    .b(__delay_data_2139__delay_2138__delay_2137__variable_681),
    .c(_cond_data_698),
    .d(__muladd_madd_odata_699)
  );

  reg [5-1:0] __delay_data_2143__delay_2142__delay_2141____variable_682;
  reg [5-1:0] __delay_data_2144__delay_2143__delay_2142____variable_682;
  reg [5-1:0] __delay_data_2145__delay_2144__delay_2143____variable_682;
  reg [5-1:0] __delay_data_2146__delay_2145__delay_2144____variable_682;
  reg signed [32-1:0] _sra_data_700;
  wire signed [32-1:0] mul_32_z_data;
  assign mul_32_z_data = _sra_data_700;
  wire signed [16-1:0] mul_33_x_data;
  wire signed [16-1:0] mul_33_y_data;
  wire [5-1:0] mul_33_rshift_data;
  reg __mul_33_stream_ivalid_1;
  reg __mul_33_stream_ivalid_2;
  reg __mul_33_stream_ivalid_3;
  reg __mul_33_stream_ivalid_4;
  reg __mul_33_stream_ivalid_5;
  reg __mul_33_stream_ivalid_6;
  reg __mul_33_stream_ivalid_7;
  reg __mul_33_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_704;
  reg [5-1:0] _minus_data_706;
  reg [1-1:0] _greatereq_data_717;
  reg signed [16-1:0] __delay_data_2153__variable_701;
  reg signed [16-1:0] __delay_data_2156__variable_702;
  reg [5-1:0] __delay_data_2159__variable_703;
  reg signed [34-1:0] _sll_data_708;
  reg [1-1:0] __delay_data_2150_greaterthan_704;
  reg [1-1:0] __delay_data_2151_greatereq_717;
  reg signed [16-1:0] __delay_data_2154__delay_2153__variable_701;
  reg signed [16-1:0] __delay_data_2157__delay_2156__variable_702;
  reg [5-1:0] __delay_data_2160__delay_2159__variable_703;
  reg signed [32-1:0] _cond_data_714;
  reg [1-1:0] __delay_data_2152__delay_2151_greatereq_717;
  reg signed [16-1:0] __delay_data_2155__delay_2154__delay_2153__variable_701;
  reg signed [16-1:0] __delay_data_2158__delay_2157__delay_2156__variable_702;
  reg [5-1:0] __delay_data_2161__delay_2160__delay_2159__variable_703;
  wire signed [16-1:0] _uminus_data_716;
  assign _uminus_data_716 = -_cond_data_714;
  wire signed [16-1:0] _cond_data_719;
  assign _cond_data_719 = (__delay_data_2152__delay_2151_greatereq_717)? _cond_data_714 : _uminus_data_716;
  wire signed [32-1:0] __muladd_madd_odata_720;
  reg signed [32-1:0] __muladd_madd_odata_reg_720;
  wire signed [32-1:0] __muladd_data_720;
  assign __muladd_data_720 = __muladd_madd_odata_reg_720;
  wire __muladd_madd_update_720;
  assign __muladd_madd_update_720 = _mul_33_stream_oready;

  madd_25
  __muladd_madd_720
  (
    .CLK(CLK),
    .update(__muladd_madd_update_720),
    .a(__delay_data_2155__delay_2154__delay_2153__variable_701),
    .b(__delay_data_2158__delay_2157__delay_2156__variable_702),
    .c(_cond_data_719),
    .d(__muladd_madd_odata_720)
  );

  reg [5-1:0] __delay_data_2162__delay_2161__delay_2160____variable_703;
  reg [5-1:0] __delay_data_2163__delay_2162__delay_2161____variable_703;
  reg [5-1:0] __delay_data_2164__delay_2163__delay_2162____variable_703;
  reg [5-1:0] __delay_data_2165__delay_2164__delay_2163____variable_703;
  reg signed [32-1:0] _sra_data_721;
  wire signed [32-1:0] mul_33_z_data;
  assign mul_33_z_data = _sra_data_721;
  wire signed [16-1:0] mul_34_x_data;
  wire signed [16-1:0] mul_34_y_data;
  wire [5-1:0] mul_34_rshift_data;
  reg __mul_34_stream_ivalid_1;
  reg __mul_34_stream_ivalid_2;
  reg __mul_34_stream_ivalid_3;
  reg __mul_34_stream_ivalid_4;
  reg __mul_34_stream_ivalid_5;
  reg __mul_34_stream_ivalid_6;
  reg __mul_34_stream_ivalid_7;
  reg __mul_34_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_725;
  reg [5-1:0] _minus_data_727;
  reg [1-1:0] _greatereq_data_738;
  reg signed [16-1:0] __delay_data_2172__variable_722;
  reg signed [16-1:0] __delay_data_2175__variable_723;
  reg [5-1:0] __delay_data_2178__variable_724;
  reg signed [34-1:0] _sll_data_729;
  reg [1-1:0] __delay_data_2169_greaterthan_725;
  reg [1-1:0] __delay_data_2170_greatereq_738;
  reg signed [16-1:0] __delay_data_2173__delay_2172__variable_722;
  reg signed [16-1:0] __delay_data_2176__delay_2175__variable_723;
  reg [5-1:0] __delay_data_2179__delay_2178__variable_724;
  reg signed [32-1:0] _cond_data_735;
  reg [1-1:0] __delay_data_2171__delay_2170_greatereq_738;
  reg signed [16-1:0] __delay_data_2174__delay_2173__delay_2172__variable_722;
  reg signed [16-1:0] __delay_data_2177__delay_2176__delay_2175__variable_723;
  reg [5-1:0] __delay_data_2180__delay_2179__delay_2178__variable_724;
  wire signed [16-1:0] _uminus_data_737;
  assign _uminus_data_737 = -_cond_data_735;
  wire signed [16-1:0] _cond_data_740;
  assign _cond_data_740 = (__delay_data_2171__delay_2170_greatereq_738)? _cond_data_735 : _uminus_data_737;
  wire signed [32-1:0] __muladd_madd_odata_741;
  reg signed [32-1:0] __muladd_madd_odata_reg_741;
  wire signed [32-1:0] __muladd_data_741;
  assign __muladd_data_741 = __muladd_madd_odata_reg_741;
  wire __muladd_madd_update_741;
  assign __muladd_madd_update_741 = _mul_34_stream_oready;

  madd_26
  __muladd_madd_741
  (
    .CLK(CLK),
    .update(__muladd_madd_update_741),
    .a(__delay_data_2174__delay_2173__delay_2172__variable_722),
    .b(__delay_data_2177__delay_2176__delay_2175__variable_723),
    .c(_cond_data_740),
    .d(__muladd_madd_odata_741)
  );

  reg [5-1:0] __delay_data_2181__delay_2180__delay_2179____variable_724;
  reg [5-1:0] __delay_data_2182__delay_2181__delay_2180____variable_724;
  reg [5-1:0] __delay_data_2183__delay_2182__delay_2181____variable_724;
  reg [5-1:0] __delay_data_2184__delay_2183__delay_2182____variable_724;
  reg signed [32-1:0] _sra_data_742;
  wire signed [32-1:0] mul_34_z_data;
  assign mul_34_z_data = _sra_data_742;
  wire signed [16-1:0] mul_35_x_data;
  wire signed [16-1:0] mul_35_y_data;
  wire [5-1:0] mul_35_rshift_data;
  reg __mul_35_stream_ivalid_1;
  reg __mul_35_stream_ivalid_2;
  reg __mul_35_stream_ivalid_3;
  reg __mul_35_stream_ivalid_4;
  reg __mul_35_stream_ivalid_5;
  reg __mul_35_stream_ivalid_6;
  reg __mul_35_stream_ivalid_7;
  reg __mul_35_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_746;
  reg [5-1:0] _minus_data_748;
  reg [1-1:0] _greatereq_data_759;
  reg signed [16-1:0] __delay_data_2209__variable_743;
  reg signed [16-1:0] __delay_data_2212__variable_744;
  reg [5-1:0] __delay_data_2215__variable_745;
  reg signed [34-1:0] _sll_data_750;
  reg [1-1:0] __delay_data_2206_greaterthan_746;
  reg [1-1:0] __delay_data_2207_greatereq_759;
  reg signed [16-1:0] __delay_data_2210__delay_2209__variable_743;
  reg signed [16-1:0] __delay_data_2213__delay_2212__variable_744;
  reg [5-1:0] __delay_data_2216__delay_2215__variable_745;
  reg signed [32-1:0] _cond_data_756;
  reg [1-1:0] __delay_data_2208__delay_2207_greatereq_759;
  reg signed [16-1:0] __delay_data_2211__delay_2210__delay_2209__variable_743;
  reg signed [16-1:0] __delay_data_2214__delay_2213__delay_2212__variable_744;
  reg [5-1:0] __delay_data_2217__delay_2216__delay_2215__variable_745;
  wire signed [16-1:0] _uminus_data_758;
  assign _uminus_data_758 = -_cond_data_756;
  wire signed [16-1:0] _cond_data_761;
  assign _cond_data_761 = (__delay_data_2208__delay_2207_greatereq_759)? _cond_data_756 : _uminus_data_758;
  wire signed [32-1:0] __muladd_madd_odata_762;
  reg signed [32-1:0] __muladd_madd_odata_reg_762;
  wire signed [32-1:0] __muladd_data_762;
  assign __muladd_data_762 = __muladd_madd_odata_reg_762;
  wire __muladd_madd_update_762;
  assign __muladd_madd_update_762 = _mul_35_stream_oready;

  madd_27
  __muladd_madd_762
  (
    .CLK(CLK),
    .update(__muladd_madd_update_762),
    .a(__delay_data_2211__delay_2210__delay_2209__variable_743),
    .b(__delay_data_2214__delay_2213__delay_2212__variable_744),
    .c(_cond_data_761),
    .d(__muladd_madd_odata_762)
  );

  reg [5-1:0] __delay_data_2218__delay_2217__delay_2216____variable_745;
  reg [5-1:0] __delay_data_2219__delay_2218__delay_2217____variable_745;
  reg [5-1:0] __delay_data_2220__delay_2219__delay_2218____variable_745;
  reg [5-1:0] __delay_data_2221__delay_2220__delay_2219____variable_745;
  reg signed [32-1:0] _sra_data_763;
  wire signed [32-1:0] mul_35_z_data;
  assign mul_35_z_data = _sra_data_763;
  wire signed [16-1:0] mul_36_x_data;
  wire signed [16-1:0] mul_36_y_data;
  wire [5-1:0] mul_36_rshift_data;
  reg __mul_36_stream_ivalid_1;
  reg __mul_36_stream_ivalid_2;
  reg __mul_36_stream_ivalid_3;
  reg __mul_36_stream_ivalid_4;
  reg __mul_36_stream_ivalid_5;
  reg __mul_36_stream_ivalid_6;
  reg __mul_36_stream_ivalid_7;
  reg __mul_36_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_767;
  reg [5-1:0] _minus_data_769;
  reg [1-1:0] _greatereq_data_780;
  reg signed [16-1:0] __delay_data_2228__variable_764;
  reg signed [16-1:0] __delay_data_2231__variable_765;
  reg [5-1:0] __delay_data_2234__variable_766;
  reg signed [34-1:0] _sll_data_771;
  reg [1-1:0] __delay_data_2225_greaterthan_767;
  reg [1-1:0] __delay_data_2226_greatereq_780;
  reg signed [16-1:0] __delay_data_2229__delay_2228__variable_764;
  reg signed [16-1:0] __delay_data_2232__delay_2231__variable_765;
  reg [5-1:0] __delay_data_2235__delay_2234__variable_766;
  reg signed [32-1:0] _cond_data_777;
  reg [1-1:0] __delay_data_2227__delay_2226_greatereq_780;
  reg signed [16-1:0] __delay_data_2230__delay_2229__delay_2228__variable_764;
  reg signed [16-1:0] __delay_data_2233__delay_2232__delay_2231__variable_765;
  reg [5-1:0] __delay_data_2236__delay_2235__delay_2234__variable_766;
  wire signed [16-1:0] _uminus_data_779;
  assign _uminus_data_779 = -_cond_data_777;
  wire signed [16-1:0] _cond_data_782;
  assign _cond_data_782 = (__delay_data_2227__delay_2226_greatereq_780)? _cond_data_777 : _uminus_data_779;
  wire signed [32-1:0] __muladd_madd_odata_783;
  reg signed [32-1:0] __muladd_madd_odata_reg_783;
  wire signed [32-1:0] __muladd_data_783;
  assign __muladd_data_783 = __muladd_madd_odata_reg_783;
  wire __muladd_madd_update_783;
  assign __muladd_madd_update_783 = _mul_36_stream_oready;

  madd_28
  __muladd_madd_783
  (
    .CLK(CLK),
    .update(__muladd_madd_update_783),
    .a(__delay_data_2230__delay_2229__delay_2228__variable_764),
    .b(__delay_data_2233__delay_2232__delay_2231__variable_765),
    .c(_cond_data_782),
    .d(__muladd_madd_odata_783)
  );

  reg [5-1:0] __delay_data_2237__delay_2236__delay_2235____variable_766;
  reg [5-1:0] __delay_data_2238__delay_2237__delay_2236____variable_766;
  reg [5-1:0] __delay_data_2239__delay_2238__delay_2237____variable_766;
  reg [5-1:0] __delay_data_2240__delay_2239__delay_2238____variable_766;
  reg signed [32-1:0] _sra_data_784;
  wire signed [32-1:0] mul_36_z_data;
  assign mul_36_z_data = _sra_data_784;
  wire signed [16-1:0] mul_37_x_data;
  wire signed [16-1:0] mul_37_y_data;
  wire [5-1:0] mul_37_rshift_data;
  reg __mul_37_stream_ivalid_1;
  reg __mul_37_stream_ivalid_2;
  reg __mul_37_stream_ivalid_3;
  reg __mul_37_stream_ivalid_4;
  reg __mul_37_stream_ivalid_5;
  reg __mul_37_stream_ivalid_6;
  reg __mul_37_stream_ivalid_7;
  reg __mul_37_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_788;
  reg [5-1:0] _minus_data_790;
  reg [1-1:0] _greatereq_data_801;
  reg signed [16-1:0] __delay_data_2247__variable_785;
  reg signed [16-1:0] __delay_data_2250__variable_786;
  reg [5-1:0] __delay_data_2253__variable_787;
  reg signed [34-1:0] _sll_data_792;
  reg [1-1:0] __delay_data_2244_greaterthan_788;
  reg [1-1:0] __delay_data_2245_greatereq_801;
  reg signed [16-1:0] __delay_data_2248__delay_2247__variable_785;
  reg signed [16-1:0] __delay_data_2251__delay_2250__variable_786;
  reg [5-1:0] __delay_data_2254__delay_2253__variable_787;
  reg signed [32-1:0] _cond_data_798;
  reg [1-1:0] __delay_data_2246__delay_2245_greatereq_801;
  reg signed [16-1:0] __delay_data_2249__delay_2248__delay_2247__variable_785;
  reg signed [16-1:0] __delay_data_2252__delay_2251__delay_2250__variable_786;
  reg [5-1:0] __delay_data_2255__delay_2254__delay_2253__variable_787;
  wire signed [16-1:0] _uminus_data_800;
  assign _uminus_data_800 = -_cond_data_798;
  wire signed [16-1:0] _cond_data_803;
  assign _cond_data_803 = (__delay_data_2246__delay_2245_greatereq_801)? _cond_data_798 : _uminus_data_800;
  wire signed [32-1:0] __muladd_madd_odata_804;
  reg signed [32-1:0] __muladd_madd_odata_reg_804;
  wire signed [32-1:0] __muladd_data_804;
  assign __muladd_data_804 = __muladd_madd_odata_reg_804;
  wire __muladd_madd_update_804;
  assign __muladd_madd_update_804 = _mul_37_stream_oready;

  madd_29
  __muladd_madd_804
  (
    .CLK(CLK),
    .update(__muladd_madd_update_804),
    .a(__delay_data_2249__delay_2248__delay_2247__variable_785),
    .b(__delay_data_2252__delay_2251__delay_2250__variable_786),
    .c(_cond_data_803),
    .d(__muladd_madd_odata_804)
  );

  reg [5-1:0] __delay_data_2256__delay_2255__delay_2254____variable_787;
  reg [5-1:0] __delay_data_2257__delay_2256__delay_2255____variable_787;
  reg [5-1:0] __delay_data_2258__delay_2257__delay_2256____variable_787;
  reg [5-1:0] __delay_data_2259__delay_2258__delay_2257____variable_787;
  reg signed [32-1:0] _sra_data_805;
  wire signed [32-1:0] mul_37_z_data;
  assign mul_37_z_data = _sra_data_805;
  wire signed [16-1:0] mul_38_x_data;
  wire signed [16-1:0] mul_38_y_data;
  wire [5-1:0] mul_38_rshift_data;
  reg __mul_38_stream_ivalid_1;
  reg __mul_38_stream_ivalid_2;
  reg __mul_38_stream_ivalid_3;
  reg __mul_38_stream_ivalid_4;
  reg __mul_38_stream_ivalid_5;
  reg __mul_38_stream_ivalid_6;
  reg __mul_38_stream_ivalid_7;
  reg __mul_38_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_809;
  reg [5-1:0] _minus_data_811;
  reg [1-1:0] _greatereq_data_822;
  reg signed [16-1:0] __delay_data_2266__variable_806;
  reg signed [16-1:0] __delay_data_2269__variable_807;
  reg [5-1:0] __delay_data_2272__variable_808;
  reg signed [34-1:0] _sll_data_813;
  reg [1-1:0] __delay_data_2263_greaterthan_809;
  reg [1-1:0] __delay_data_2264_greatereq_822;
  reg signed [16-1:0] __delay_data_2267__delay_2266__variable_806;
  reg signed [16-1:0] __delay_data_2270__delay_2269__variable_807;
  reg [5-1:0] __delay_data_2273__delay_2272__variable_808;
  reg signed [32-1:0] _cond_data_819;
  reg [1-1:0] __delay_data_2265__delay_2264_greatereq_822;
  reg signed [16-1:0] __delay_data_2268__delay_2267__delay_2266__variable_806;
  reg signed [16-1:0] __delay_data_2271__delay_2270__delay_2269__variable_807;
  reg [5-1:0] __delay_data_2274__delay_2273__delay_2272__variable_808;
  wire signed [16-1:0] _uminus_data_821;
  assign _uminus_data_821 = -_cond_data_819;
  wire signed [16-1:0] _cond_data_824;
  assign _cond_data_824 = (__delay_data_2265__delay_2264_greatereq_822)? _cond_data_819 : _uminus_data_821;
  wire signed [32-1:0] __muladd_madd_odata_825;
  reg signed [32-1:0] __muladd_madd_odata_reg_825;
  wire signed [32-1:0] __muladd_data_825;
  assign __muladd_data_825 = __muladd_madd_odata_reg_825;
  wire __muladd_madd_update_825;
  assign __muladd_madd_update_825 = _mul_38_stream_oready;

  madd_30
  __muladd_madd_825
  (
    .CLK(CLK),
    .update(__muladd_madd_update_825),
    .a(__delay_data_2268__delay_2267__delay_2266__variable_806),
    .b(__delay_data_2271__delay_2270__delay_2269__variable_807),
    .c(_cond_data_824),
    .d(__muladd_madd_odata_825)
  );

  reg [5-1:0] __delay_data_2275__delay_2274__delay_2273____variable_808;
  reg [5-1:0] __delay_data_2276__delay_2275__delay_2274____variable_808;
  reg [5-1:0] __delay_data_2277__delay_2276__delay_2275____variable_808;
  reg [5-1:0] __delay_data_2278__delay_2277__delay_2276____variable_808;
  reg signed [32-1:0] _sra_data_826;
  wire signed [32-1:0] mul_38_z_data;
  assign mul_38_z_data = _sra_data_826;
  wire signed [16-1:0] mul_39_x_data;
  wire signed [16-1:0] mul_39_y_data;
  wire [5-1:0] mul_39_rshift_data;
  reg __mul_39_stream_ivalid_1;
  reg __mul_39_stream_ivalid_2;
  reg __mul_39_stream_ivalid_3;
  reg __mul_39_stream_ivalid_4;
  reg __mul_39_stream_ivalid_5;
  reg __mul_39_stream_ivalid_6;
  reg __mul_39_stream_ivalid_7;
  reg __mul_39_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_830;
  reg [5-1:0] _minus_data_832;
  reg [1-1:0] _greatereq_data_843;
  reg signed [16-1:0] __delay_data_2285__variable_827;
  reg signed [16-1:0] __delay_data_2288__variable_828;
  reg [5-1:0] __delay_data_2291__variable_829;
  reg signed [34-1:0] _sll_data_834;
  reg [1-1:0] __delay_data_2282_greaterthan_830;
  reg [1-1:0] __delay_data_2283_greatereq_843;
  reg signed [16-1:0] __delay_data_2286__delay_2285__variable_827;
  reg signed [16-1:0] __delay_data_2289__delay_2288__variable_828;
  reg [5-1:0] __delay_data_2292__delay_2291__variable_829;
  reg signed [32-1:0] _cond_data_840;
  reg [1-1:0] __delay_data_2284__delay_2283_greatereq_843;
  reg signed [16-1:0] __delay_data_2287__delay_2286__delay_2285__variable_827;
  reg signed [16-1:0] __delay_data_2290__delay_2289__delay_2288__variable_828;
  reg [5-1:0] __delay_data_2293__delay_2292__delay_2291__variable_829;
  wire signed [16-1:0] _uminus_data_842;
  assign _uminus_data_842 = -_cond_data_840;
  wire signed [16-1:0] _cond_data_845;
  assign _cond_data_845 = (__delay_data_2284__delay_2283_greatereq_843)? _cond_data_840 : _uminus_data_842;
  wire signed [32-1:0] __muladd_madd_odata_846;
  reg signed [32-1:0] __muladd_madd_odata_reg_846;
  wire signed [32-1:0] __muladd_data_846;
  assign __muladd_data_846 = __muladd_madd_odata_reg_846;
  wire __muladd_madd_update_846;
  assign __muladd_madd_update_846 = _mul_39_stream_oready;

  madd_31
  __muladd_madd_846
  (
    .CLK(CLK),
    .update(__muladd_madd_update_846),
    .a(__delay_data_2287__delay_2286__delay_2285__variable_827),
    .b(__delay_data_2290__delay_2289__delay_2288__variable_828),
    .c(_cond_data_845),
    .d(__muladd_madd_odata_846)
  );

  reg [5-1:0] __delay_data_2294__delay_2293__delay_2292____variable_829;
  reg [5-1:0] __delay_data_2295__delay_2294__delay_2293____variable_829;
  reg [5-1:0] __delay_data_2296__delay_2295__delay_2294____variable_829;
  reg [5-1:0] __delay_data_2297__delay_2296__delay_2295____variable_829;
  reg signed [32-1:0] _sra_data_847;
  wire signed [32-1:0] mul_39_z_data;
  assign mul_39_z_data = _sra_data_847;
  wire signed [16-1:0] mul_40_x_data;
  wire signed [16-1:0] mul_40_y_data;
  wire [5-1:0] mul_40_rshift_data;
  reg __mul_40_stream_ivalid_1;
  reg __mul_40_stream_ivalid_2;
  reg __mul_40_stream_ivalid_3;
  reg __mul_40_stream_ivalid_4;
  reg __mul_40_stream_ivalid_5;
  reg __mul_40_stream_ivalid_6;
  reg __mul_40_stream_ivalid_7;
  reg __mul_40_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_851;
  reg [5-1:0] _minus_data_853;
  reg [1-1:0] _greatereq_data_864;
  reg signed [16-1:0] __delay_data_2304__variable_848;
  reg signed [16-1:0] __delay_data_2307__variable_849;
  reg [5-1:0] __delay_data_2310__variable_850;
  reg signed [34-1:0] _sll_data_855;
  reg [1-1:0] __delay_data_2301_greaterthan_851;
  reg [1-1:0] __delay_data_2302_greatereq_864;
  reg signed [16-1:0] __delay_data_2305__delay_2304__variable_848;
  reg signed [16-1:0] __delay_data_2308__delay_2307__variable_849;
  reg [5-1:0] __delay_data_2311__delay_2310__variable_850;
  reg signed [32-1:0] _cond_data_861;
  reg [1-1:0] __delay_data_2303__delay_2302_greatereq_864;
  reg signed [16-1:0] __delay_data_2306__delay_2305__delay_2304__variable_848;
  reg signed [16-1:0] __delay_data_2309__delay_2308__delay_2307__variable_849;
  reg [5-1:0] __delay_data_2312__delay_2311__delay_2310__variable_850;
  wire signed [16-1:0] _uminus_data_863;
  assign _uminus_data_863 = -_cond_data_861;
  wire signed [16-1:0] _cond_data_866;
  assign _cond_data_866 = (__delay_data_2303__delay_2302_greatereq_864)? _cond_data_861 : _uminus_data_863;
  wire signed [32-1:0] __muladd_madd_odata_867;
  reg signed [32-1:0] __muladd_madd_odata_reg_867;
  wire signed [32-1:0] __muladd_data_867;
  assign __muladd_data_867 = __muladd_madd_odata_reg_867;
  wire __muladd_madd_update_867;
  assign __muladd_madd_update_867 = _mul_40_stream_oready;

  madd_32
  __muladd_madd_867
  (
    .CLK(CLK),
    .update(__muladd_madd_update_867),
    .a(__delay_data_2306__delay_2305__delay_2304__variable_848),
    .b(__delay_data_2309__delay_2308__delay_2307__variable_849),
    .c(_cond_data_866),
    .d(__muladd_madd_odata_867)
  );

  reg [5-1:0] __delay_data_2313__delay_2312__delay_2311____variable_850;
  reg [5-1:0] __delay_data_2314__delay_2313__delay_2312____variable_850;
  reg [5-1:0] __delay_data_2315__delay_2314__delay_2313____variable_850;
  reg [5-1:0] __delay_data_2316__delay_2315__delay_2314____variable_850;
  reg signed [32-1:0] _sra_data_868;
  wire signed [32-1:0] mul_40_z_data;
  assign mul_40_z_data = _sra_data_868;
  wire signed [16-1:0] mul_41_x_data;
  wire signed [16-1:0] mul_41_y_data;
  wire [5-1:0] mul_41_rshift_data;
  reg __mul_41_stream_ivalid_1;
  reg __mul_41_stream_ivalid_2;
  reg __mul_41_stream_ivalid_3;
  reg __mul_41_stream_ivalid_4;
  reg __mul_41_stream_ivalid_5;
  reg __mul_41_stream_ivalid_6;
  reg __mul_41_stream_ivalid_7;
  reg __mul_41_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_872;
  reg [5-1:0] _minus_data_874;
  reg [1-1:0] _greatereq_data_885;
  reg signed [16-1:0] __delay_data_2323__variable_869;
  reg signed [16-1:0] __delay_data_2326__variable_870;
  reg [5-1:0] __delay_data_2329__variable_871;
  reg signed [34-1:0] _sll_data_876;
  reg [1-1:0] __delay_data_2320_greaterthan_872;
  reg [1-1:0] __delay_data_2321_greatereq_885;
  reg signed [16-1:0] __delay_data_2324__delay_2323__variable_869;
  reg signed [16-1:0] __delay_data_2327__delay_2326__variable_870;
  reg [5-1:0] __delay_data_2330__delay_2329__variable_871;
  reg signed [32-1:0] _cond_data_882;
  reg [1-1:0] __delay_data_2322__delay_2321_greatereq_885;
  reg signed [16-1:0] __delay_data_2325__delay_2324__delay_2323__variable_869;
  reg signed [16-1:0] __delay_data_2328__delay_2327__delay_2326__variable_870;
  reg [5-1:0] __delay_data_2331__delay_2330__delay_2329__variable_871;
  wire signed [16-1:0] _uminus_data_884;
  assign _uminus_data_884 = -_cond_data_882;
  wire signed [16-1:0] _cond_data_887;
  assign _cond_data_887 = (__delay_data_2322__delay_2321_greatereq_885)? _cond_data_882 : _uminus_data_884;
  wire signed [32-1:0] __muladd_madd_odata_888;
  reg signed [32-1:0] __muladd_madd_odata_reg_888;
  wire signed [32-1:0] __muladd_data_888;
  assign __muladd_data_888 = __muladd_madd_odata_reg_888;
  wire __muladd_madd_update_888;
  assign __muladd_madd_update_888 = _mul_41_stream_oready;

  madd_33
  __muladd_madd_888
  (
    .CLK(CLK),
    .update(__muladd_madd_update_888),
    .a(__delay_data_2325__delay_2324__delay_2323__variable_869),
    .b(__delay_data_2328__delay_2327__delay_2326__variable_870),
    .c(_cond_data_887),
    .d(__muladd_madd_odata_888)
  );

  reg [5-1:0] __delay_data_2332__delay_2331__delay_2330____variable_871;
  reg [5-1:0] __delay_data_2333__delay_2332__delay_2331____variable_871;
  reg [5-1:0] __delay_data_2334__delay_2333__delay_2332____variable_871;
  reg [5-1:0] __delay_data_2335__delay_2334__delay_2333____variable_871;
  reg signed [32-1:0] _sra_data_889;
  wire signed [32-1:0] mul_41_z_data;
  assign mul_41_z_data = _sra_data_889;
  wire signed [16-1:0] mul_42_x_data;
  wire signed [16-1:0] mul_42_y_data;
  wire [5-1:0] mul_42_rshift_data;
  reg __mul_42_stream_ivalid_1;
  reg __mul_42_stream_ivalid_2;
  reg __mul_42_stream_ivalid_3;
  reg __mul_42_stream_ivalid_4;
  reg __mul_42_stream_ivalid_5;
  reg __mul_42_stream_ivalid_6;
  reg __mul_42_stream_ivalid_7;
  reg __mul_42_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_893;
  reg [5-1:0] _minus_data_895;
  reg [1-1:0] _greatereq_data_906;
  reg signed [16-1:0] __delay_data_2342__variable_890;
  reg signed [16-1:0] __delay_data_2345__variable_891;
  reg [5-1:0] __delay_data_2348__variable_892;
  reg signed [34-1:0] _sll_data_897;
  reg [1-1:0] __delay_data_2339_greaterthan_893;
  reg [1-1:0] __delay_data_2340_greatereq_906;
  reg signed [16-1:0] __delay_data_2343__delay_2342__variable_890;
  reg signed [16-1:0] __delay_data_2346__delay_2345__variable_891;
  reg [5-1:0] __delay_data_2349__delay_2348__variable_892;
  reg signed [32-1:0] _cond_data_903;
  reg [1-1:0] __delay_data_2341__delay_2340_greatereq_906;
  reg signed [16-1:0] __delay_data_2344__delay_2343__delay_2342__variable_890;
  reg signed [16-1:0] __delay_data_2347__delay_2346__delay_2345__variable_891;
  reg [5-1:0] __delay_data_2350__delay_2349__delay_2348__variable_892;
  wire signed [16-1:0] _uminus_data_905;
  assign _uminus_data_905 = -_cond_data_903;
  wire signed [16-1:0] _cond_data_908;
  assign _cond_data_908 = (__delay_data_2341__delay_2340_greatereq_906)? _cond_data_903 : _uminus_data_905;
  wire signed [32-1:0] __muladd_madd_odata_909;
  reg signed [32-1:0] __muladd_madd_odata_reg_909;
  wire signed [32-1:0] __muladd_data_909;
  assign __muladd_data_909 = __muladd_madd_odata_reg_909;
  wire __muladd_madd_update_909;
  assign __muladd_madd_update_909 = _mul_42_stream_oready;

  madd_34
  __muladd_madd_909
  (
    .CLK(CLK),
    .update(__muladd_madd_update_909),
    .a(__delay_data_2344__delay_2343__delay_2342__variable_890),
    .b(__delay_data_2347__delay_2346__delay_2345__variable_891),
    .c(_cond_data_908),
    .d(__muladd_madd_odata_909)
  );

  reg [5-1:0] __delay_data_2351__delay_2350__delay_2349____variable_892;
  reg [5-1:0] __delay_data_2352__delay_2351__delay_2350____variable_892;
  reg [5-1:0] __delay_data_2353__delay_2352__delay_2351____variable_892;
  reg [5-1:0] __delay_data_2354__delay_2353__delay_2352____variable_892;
  reg signed [32-1:0] _sra_data_910;
  wire signed [32-1:0] mul_42_z_data;
  assign mul_42_z_data = _sra_data_910;
  wire signed [16-1:0] mul_43_x_data;
  wire signed [16-1:0] mul_43_y_data;
  wire [5-1:0] mul_43_rshift_data;
  reg __mul_43_stream_ivalid_1;
  reg __mul_43_stream_ivalid_2;
  reg __mul_43_stream_ivalid_3;
  reg __mul_43_stream_ivalid_4;
  reg __mul_43_stream_ivalid_5;
  reg __mul_43_stream_ivalid_6;
  reg __mul_43_stream_ivalid_7;
  reg __mul_43_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_914;
  reg [5-1:0] _minus_data_916;
  reg [1-1:0] _greatereq_data_927;
  reg signed [16-1:0] __delay_data_2361__variable_911;
  reg signed [16-1:0] __delay_data_2364__variable_912;
  reg [5-1:0] __delay_data_2367__variable_913;
  reg signed [34-1:0] _sll_data_918;
  reg [1-1:0] __delay_data_2358_greaterthan_914;
  reg [1-1:0] __delay_data_2359_greatereq_927;
  reg signed [16-1:0] __delay_data_2362__delay_2361__variable_911;
  reg signed [16-1:0] __delay_data_2365__delay_2364__variable_912;
  reg [5-1:0] __delay_data_2368__delay_2367__variable_913;
  reg signed [32-1:0] _cond_data_924;
  reg [1-1:0] __delay_data_2360__delay_2359_greatereq_927;
  reg signed [16-1:0] __delay_data_2363__delay_2362__delay_2361__variable_911;
  reg signed [16-1:0] __delay_data_2366__delay_2365__delay_2364__variable_912;
  reg [5-1:0] __delay_data_2369__delay_2368__delay_2367__variable_913;
  wire signed [16-1:0] _uminus_data_926;
  assign _uminus_data_926 = -_cond_data_924;
  wire signed [16-1:0] _cond_data_929;
  assign _cond_data_929 = (__delay_data_2360__delay_2359_greatereq_927)? _cond_data_924 : _uminus_data_926;
  wire signed [32-1:0] __muladd_madd_odata_930;
  reg signed [32-1:0] __muladd_madd_odata_reg_930;
  wire signed [32-1:0] __muladd_data_930;
  assign __muladd_data_930 = __muladd_madd_odata_reg_930;
  wire __muladd_madd_update_930;
  assign __muladd_madd_update_930 = _mul_43_stream_oready;

  madd_35
  __muladd_madd_930
  (
    .CLK(CLK),
    .update(__muladd_madd_update_930),
    .a(__delay_data_2363__delay_2362__delay_2361__variable_911),
    .b(__delay_data_2366__delay_2365__delay_2364__variable_912),
    .c(_cond_data_929),
    .d(__muladd_madd_odata_930)
  );

  reg [5-1:0] __delay_data_2370__delay_2369__delay_2368____variable_913;
  reg [5-1:0] __delay_data_2371__delay_2370__delay_2369____variable_913;
  reg [5-1:0] __delay_data_2372__delay_2371__delay_2370____variable_913;
  reg [5-1:0] __delay_data_2373__delay_2372__delay_2371____variable_913;
  reg signed [32-1:0] _sra_data_931;
  wire signed [32-1:0] mul_43_z_data;
  assign mul_43_z_data = _sra_data_931;
  wire signed [64-1:0] add_tree_5_var0_data;
  wire signed [64-1:0] add_tree_5_var1_data;
  wire signed [64-1:0] add_tree_5_var2_data;
  wire signed [64-1:0] add_tree_5_var3_data;
  wire signed [64-1:0] add_tree_5_var4_data;
  wire signed [64-1:0] add_tree_5_var5_data;
  wire signed [64-1:0] add_tree_5_var6_data;
  wire signed [64-1:0] add_tree_5_var7_data;
  wire signed [64-1:0] add_tree_5_var8_data;
  wire signed [64-1:0] add_tree_5_var9_data;
  wire signed [64-1:0] add_tree_5_var10_data;
  wire signed [64-1:0] add_tree_5_var11_data;
  wire signed [64-1:0] add_tree_5_var12_data;
  wire signed [64-1:0] add_tree_5_var13_data;
  wire signed [64-1:0] add_tree_5_var14_data;
  wire signed [64-1:0] add_tree_5_var15_data;
  wire signed [64-1:0] add_tree_5_var16_data;
  wire signed [64-1:0] add_tree_5_var17_data;
  reg __add_tree_5_stream_ivalid_1;
  reg __add_tree_5_stream_ivalid_2;
  reg __add_tree_5_stream_ivalid_3;
  reg signed [64-1:0] __plusn_data_99;
  reg signed [64-1:0] __plusn_data_100;
  reg signed [64-1:0] __plusn_data_101;
  reg signed [64-1:0] __plusn_data_103;
  reg signed [64-1:0] __plusn_data_104;
  reg signed [64-1:0] __plusn_data_105;
  reg signed [64-1:0] __plusn_data_102;
  reg signed [64-1:0] __plusn_data_106;
  reg signed [64-1:0] __plusn_data_107;
  wire signed [64-1:0] add_tree_5_sum_data;
  assign add_tree_5_sum_data = __plusn_data_107;
  wire signed [64-1:0] acc_1_x_data;
  wire [7-1:0] acc_1_rshift_data;
  wire [32-1:0] acc_1_size_data;
  wire [1-1:0] acc_1__reduce_reset_data;
  reg __acc_1_stream_ivalid_1;
  reg __acc_1_stream_ivalid_2;
  reg __acc_1_stream_ivalid_3;
  reg __acc_1_stream_ivalid_4;
  reg __acc_1_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_25;
  reg [7-1:0] _minus_data_27;
  reg signed [64-1:0] _reduceadd_data_38;
  reg [33-1:0] _reduceadd_count_38;
  reg _reduceadd_prev_count_max_38;
  wire _reduceadd_reset_cond_38;
  assign _reduceadd_reset_cond_38 = acc_1__reduce_reset_data || _reduceadd_prev_count_max_38;
  wire [33-1:0] _reduceadd_current_count_38;
  assign _reduceadd_current_count_38 = (_reduceadd_reset_cond_38)? 0 : _reduceadd_count_38;
  wire signed [64-1:0] _reduceadd_current_data_38;
  assign _reduceadd_current_data_38 = (_reduceadd_reset_cond_38)? 1'sd0 : _reduceadd_data_38;
  reg [1-1:0] _pulse_data_40;
  reg [33-1:0] _pulse_count_40;
  reg _pulse_prev_count_max_40;
  wire _pulse_reset_cond_40;
  assign _pulse_reset_cond_40 = acc_1__reduce_reset_data || _pulse_prev_count_max_40;
  wire [33-1:0] _pulse_current_count_40;
  assign _pulse_current_count_40 = (_pulse_reset_cond_40)? 0 : _pulse_count_40;
  wire [1-1:0] _pulse_current_data_40;
  assign _pulse_current_data_40 = (_pulse_reset_cond_40)? 1'sd0 : _pulse_data_40;
  reg [7-1:0] __delay_data_2382__variable_23;
  reg signed [130-1:0] _sll_data_29;
  reg [1-1:0] __delay_data_2379_greaterthan_25;
  reg signed [64-1:0] __delay_data_2380_reduceadd_38;
  reg [7-1:0] __delay_data_2383__delay_2382__variable_23;
  reg [1-1:0] __delay_data_2386_pulse_40;
  reg signed [64-1:0] _cond_data_35;
  reg signed [64-1:0] __delay_data_2381__delay_2380_reduceadd_38;
  reg [7-1:0] __delay_data_2384__delay_2383__delay_2382__variable_23;
  reg [1-1:0] __delay_data_2387__delay_2386_pulse_40;
  reg signed [64-1:0] _plus_data_42;
  reg [7-1:0] __delay_data_2385__delay_2384__delay_2383____variable_23;
  reg [1-1:0] __delay_data_2388__delay_2387__delay_2386_pulse_40;
  reg signed [64-1:0] _sra_data_43;
  reg [1-1:0] __delay_data_2389__delay_2388__delay_2387__delay_2386_pulse_40;
  wire signed [64-1:0] acc_1_sum_data;
  assign acc_1_sum_data = _sra_data_43;
  wire [1-1:0] acc_1_valid_data;
  assign acc_1_valid_data = __delay_data_2389__delay_2388__delay_2387__delay_2386_pulse_40;
  wire signed [64-1:0] mul_rshift_round_clip_7_x_data;
  wire signed [16-1:0] mul_rshift_round_clip_7_y_data;
  wire [7-1:0] mul_rshift_round_clip_7_rshift_data;
  reg __mul_rshift_round_clip_7_stream_ivalid_1;
  reg __mul_rshift_round_clip_7_stream_ivalid_2;
  reg __mul_rshift_round_clip_7_stream_ivalid_3;
  reg __mul_rshift_round_clip_7_stream_ivalid_4;
  reg __mul_rshift_round_clip_7_stream_ivalid_5;
  reg __mul_rshift_round_clip_7_stream_ivalid_6;
  reg __mul_rshift_round_clip_7_stream_ivalid_7;
  reg __mul_rshift_round_clip_7_stream_ivalid_8;
  wire signed [80-1:0] _times_mul_odata_145;
  reg signed [80-1:0] _times_mul_odata_reg_145;
  wire signed [80-1:0] _times_data_145;
  assign _times_data_145 = _times_mul_odata_reg_145;
  wire _times_mul_update_145;
  assign _times_mul_update_145 = _mul_rshift_round_clip_7_stream_oready;

  multiplier_1
  _times_mul_145
  (
    .CLK(CLK),
    .update(_times_mul_update_145),
    .a(mul_rshift_round_clip_7_x_data),
    .b(mul_rshift_round_clip_7_y_data),
    .c(_times_mul_odata_145)
  );

  wire [7-1:0] _minus_data_148;
  assign _minus_data_148 = mul_rshift_round_clip_7_rshift_data - 2'sd1;
  wire signed [130-1:0] _sll_data_151;
  assign _sll_data_151 = 2'sd1 << _minus_data_148;
  wire [1-1:0] _eq_data_163;
  assign _eq_data_163 = mul_rshift_round_clip_7_rshift_data == 1'sd0;
  reg signed [130-1:0] __delay_data_2395_sll_151;
  reg [7-1:0] __delay_data_2399__variable_144;
  reg [1-1:0] __delay_data_2403_eq_163;
  reg signed [130-1:0] __delay_data_2396__delay_2395_sll_151;
  reg [7-1:0] __delay_data_2400__delay_2399__variable_144;
  reg [1-1:0] __delay_data_2404__delay_2403_eq_163;
  reg signed [130-1:0] __delay_data_2397__delay_2396__delay_2395_sll_151;
  reg [7-1:0] __delay_data_2401__delay_2400__delay_2399__variable_144;
  reg [1-1:0] __delay_data_2405__delay_2404__delay_2403_eq_163;
  reg signed [130-1:0] __delay_data_2398__delay_2397__delay_2396__delay_2395_sll_151;
  reg [7-1:0] __delay_data_2402__delay_2401__delay_2400____variable_144;
  reg [1-1:0] __delay_data_2406__delay_2405__delay_2404__delay_2403_eq_163;
  wire [1-1:0] _pointer_data_146;
  assign _pointer_data_146 = _times_data_145[8'sd79];
  wire signed [2-1:0] _cond_data_158;
  assign _cond_data_158 = (_pointer_data_146)? -2'sd1 : 1'sd0;
  wire signed [81-1:0] _plus_data_159;
  assign _plus_data_159 = _times_data_145 + __delay_data_2398__delay_2397__delay_2396__delay_2395_sll_151;
  wire signed [81-1:0] _plus_data_160;
  assign _plus_data_160 = _plus_data_159 + _cond_data_158;
  wire signed [80-1:0] _sra_data_161;
  assign _sra_data_161 = _plus_data_160 >>> __delay_data_2402__delay_2401__delay_2400____variable_144;
  reg signed [80-1:0] _cond_data_164;
  reg [1-1:0] _greaterthan_data_165;
  reg [1-1:0] _lessthan_data_169;
  reg [1-1:0] _greatereq_data_173;
  reg signed [80-1:0] __delay_data_2407_cond_164;
  reg signed [80-1:0] _cond_data_167;
  reg signed [80-1:0] _cond_data_171;
  reg [1-1:0] __delay_data_2408_greatereq_173;
  reg signed [16-1:0] _cond_data_175;
  wire signed [16-1:0] mul_rshift_round_clip_7_z_data;
  assign mul_rshift_round_clip_7_z_data = _cond_data_175;
  reg [33-1:0] _stream_conv2d_4_sink_89_sink_count;
  reg [5-1:0] _stream_conv2d_4_sink_89_sink_mode;
  reg [16-1:0] _stream_conv2d_4_sink_89_sink_generator_id;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_offset;
  reg [33-1:0] _stream_conv2d_4_sink_89_sink_size;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_stride;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_4_sink_89_sink_size_buf;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_4_sink_89_sink_sel;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_waddr;
  reg _stream_conv2d_4_sink_89_sink_wenable;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_wdata;
  reg _stream_conv2d_4_sink_89_sink_fifo_enq;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_fifo_wdata;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_immediate;
  reg [33-1:0] _stream_conv2d_4_sink_90_sink_count;
  reg [5-1:0] _stream_conv2d_4_sink_90_sink_mode;
  reg [16-1:0] _stream_conv2d_4_sink_90_sink_generator_id;
  reg [32-1:0] _stream_conv2d_4_sink_90_sink_offset;
  reg [33-1:0] _stream_conv2d_4_sink_90_sink_size;
  reg [32-1:0] _stream_conv2d_4_sink_90_sink_stride;
  reg [32-1:0] _stream_conv2d_4_sink_90_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_4_sink_90_sink_size_buf;
  reg [32-1:0] _stream_conv2d_4_sink_90_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_4_sink_90_sink_sel;
  reg [32-1:0] _stream_conv2d_4_sink_90_sink_waddr;
  reg _stream_conv2d_4_sink_90_sink_wenable;
  reg [1-1:0] _stream_conv2d_4_sink_90_sink_wdata;
  reg _stream_conv2d_4_sink_90_sink_fifo_enq;
  reg [1-1:0] _stream_conv2d_4_sink_90_sink_fifo_wdata;
  reg [1-1:0] _stream_conv2d_4_sink_90_sink_immediate;
  reg _stream_max_pool_serial_6_stream_ivalid;
  wire _stream_max_pool_serial_6_stream_oready;
  wire _stream_max_pool_serial_6_stream_internal_oready;
  assign _stream_max_pool_serial_6_stream_oready = _stream_max_pool_serial_6_stream_internal_oready;
  reg [32-1:0] _stream_max_pool_serial_6_fsm;
  localparam _stream_max_pool_serial_6_fsm_init = 0;
  wire _stream_max_pool_serial_6_run_flag;
  reg _stream_max_pool_serial_6_source_start;
  wire _stream_max_pool_serial_6_source_stop;
  reg _stream_max_pool_serial_6_source_busy;
  wire _stream_max_pool_serial_6_sink_start;
  wire _stream_max_pool_serial_6_sink_stop;
  wire _stream_max_pool_serial_6_sink_busy;
  wire _stream_max_pool_serial_6_busy;
  reg _stream_max_pool_serial_6_busy_reg;
  wire _stream_max_pool_serial_6_is_root;
  assign _stream_max_pool_serial_6_is_root = 1;
  reg [3-1:0] _stream_max_pool_serial_6_parameter_0_next_parameter_data;
  reg _stream_max_pool_serial_6_source_1_idle;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_count;
  reg [5-1:0] _stream_max_pool_serial_6_source_1_source_mode;
  reg [16-1:0] _stream_max_pool_serial_6_source_1_source_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_offset;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_size;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_stride;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_source_1_source_sel;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_ram_raddr;
  reg _stream_max_pool_serial_6_source_1_source_ram_renable;
  wire [32-1:0] _stream_max_pool_serial_6_source_1_source_ram_rdata;
  reg _stream_max_pool_serial_6_source_1_source_fifo_deq;
  wire [32-1:0] _stream_max_pool_serial_6_source_1_source_fifo_rdata;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_empty_data;
  reg [4-1:0] _stream_max_pool_serial_6_parameter_2_next_parameter_data;
  wire signed [16-1:0] _reduce_max_44_x_data;
  wire [32-1:0] _reduce_max_44_size_data;
  wire [1-1:0] _reduce_max_44__reduce_reset_data;
  reg ___reduce_max_44_stream_ivalid_1;
  reg signed [16-1:0] _reducemax_data_935;
  reg [33-1:0] _reducemax_count_935;
  reg _reducemax_prev_count_max_935;
  wire _reducemax_reset_cond_935;
  assign _reducemax_reset_cond_935 = _reduce_max_44__reduce_reset_data || _reducemax_prev_count_max_935;
  wire [33-1:0] _reducemax_current_count_935;
  assign _reducemax_current_count_935 = (_reducemax_reset_cond_935)? 0 : _reducemax_count_935;
  wire signed [16-1:0] _reducemax_current_data_935;
  assign _reducemax_current_data_935 = (_reducemax_reset_cond_935)? -17'sd32768 : _reducemax_data_935;
  reg [1-1:0] _pulse_data_937;
  reg [33-1:0] _pulse_count_937;
  reg _pulse_prev_count_max_937;
  wire _pulse_reset_cond_937;
  assign _pulse_reset_cond_937 = _reduce_max_44__reduce_reset_data || _pulse_prev_count_max_937;
  wire [33-1:0] _pulse_current_count_937;
  assign _pulse_current_count_937 = (_pulse_reset_cond_937)? 0 : _pulse_count_937;
  wire [1-1:0] _pulse_current_data_937;
  assign _pulse_current_data_937 = (_pulse_reset_cond_937)? 1'sd0 : _pulse_data_937;
  wire signed [16-1:0] _reduce_max_44_data_data;
  assign _reduce_max_44_data_data = _reducemax_data_935;
  wire [1-1:0] _reduce_max_44_valid_data;
  assign _reduce_max_44_valid_data = _pulse_data_937;
  wire signed [16-1:0] _reduce_max_45_x_data;
  wire [32-1:0] _reduce_max_45_size_data;
  wire [1-1:0] _reduce_max_45__reduce_reset_data;
  reg ___reduce_max_45_stream_ivalid_1;
  reg signed [16-1:0] _reducemax_data_942;
  reg [33-1:0] _reducemax_count_942;
  reg _reducemax_prev_count_max_942;
  wire _reducemax_reset_cond_942;
  assign _reducemax_reset_cond_942 = _reduce_max_45__reduce_reset_data || _reducemax_prev_count_max_942;
  wire [33-1:0] _reducemax_current_count_942;
  assign _reducemax_current_count_942 = (_reducemax_reset_cond_942)? 0 : _reducemax_count_942;
  wire signed [16-1:0] _reducemax_current_data_942;
  assign _reducemax_current_data_942 = (_reducemax_reset_cond_942)? -17'sd32768 : _reducemax_data_942;
  reg [1-1:0] _pulse_data_944;
  reg [33-1:0] _pulse_count_944;
  reg _pulse_prev_count_max_944;
  wire _pulse_reset_cond_944;
  assign _pulse_reset_cond_944 = _reduce_max_45__reduce_reset_data || _pulse_prev_count_max_944;
  wire [33-1:0] _pulse_current_count_944;
  assign _pulse_current_count_944 = (_pulse_reset_cond_944)? 0 : _pulse_count_944;
  wire [1-1:0] _pulse_current_data_944;
  assign _pulse_current_data_944 = (_pulse_reset_cond_944)? 1'sd0 : _pulse_data_944;
  wire signed [16-1:0] _reduce_max_45_data_data;
  assign _reduce_max_45_data_data = _reducemax_data_942;
  wire [1-1:0] _reduce_max_45_valid_data;
  assign _reduce_max_45_valid_data = _pulse_data_944;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_count;
  reg [5-1:0] _stream_max_pool_serial_6_sink_6_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_6_sink_6_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_size;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_sink_6_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_waddr;
  reg _stream_max_pool_serial_6_sink_6_sink_wenable;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_wdata;
  reg _stream_max_pool_serial_6_sink_6_sink_fifo_enq;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_fifo_wdata;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_immediate;
  reg [33-1:0] _stream_max_pool_serial_6_sink_7_sink_count;
  reg [5-1:0] _stream_max_pool_serial_6_sink_7_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_6_sink_7_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_6_sink_7_sink_size;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_sink_7_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_sink_7_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_6_sink_7_sink_waddr;
  reg _stream_max_pool_serial_6_sink_7_sink_wenable;
  reg [1-1:0] _stream_max_pool_serial_6_sink_7_sink_wdata;
  reg _stream_max_pool_serial_6_sink_7_sink_fifo_enq;
  reg [1-1:0] _stream_max_pool_serial_6_sink_7_sink_fifo_wdata;
  reg [1-1:0] _stream_max_pool_serial_6_sink_7_sink_immediate;
  reg _stream_matmul_16_stream_ivalid;
  wire _stream_matmul_16_stream_oready;
  wire _stream_matmul_16_stream_internal_oready;
  assign _stream_matmul_16_stream_oready = _stream_matmul_16_stream_internal_oready;
  reg [32-1:0] _stream_matmul_16_fsm;
  localparam _stream_matmul_16_fsm_init = 0;
  wire _stream_matmul_16_run_flag;
  reg _stream_matmul_16_source_start;
  wire _stream_matmul_16_source_stop;
  reg _stream_matmul_16_source_busy;
  wire _stream_matmul_16_sink_start;
  wire _stream_matmul_16_sink_stop;
  wire _stream_matmul_16_sink_busy;
  wire _stream_matmul_16_busy;
  reg _stream_matmul_16_busy_reg;
  wire _stream_matmul_16_is_root;
  assign _stream_matmul_16_is_root = 1;
  reg [14-1:0] _stream_matmul_16_parameter_0_next_parameter_data;
  reg [1-1:0] _stream_matmul_16_parameter_1_next_parameter_data;
  reg [1-1:0] _stream_matmul_16_parameter_2_next_parameter_data;
  reg [1-1:0] _stream_matmul_16_parameter_3_next_parameter_data;
  reg [2-1:0] _stream_matmul_16_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_matmul_16_parameter_6_next_parameter_data;
  reg _stream_matmul_16_source_7_idle;
  reg [33-1:0] _stream_matmul_16_source_7_source_count;
  reg [5-1:0] _stream_matmul_16_source_7_source_mode;
  reg [16-1:0] _stream_matmul_16_source_7_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_7_source_offset;
  reg [33-1:0] _stream_matmul_16_source_7_source_size;
  reg [32-1:0] _stream_matmul_16_source_7_source_stride;
  reg [32-1:0] _stream_matmul_16_source_7_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_7_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_7_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_7_source_sel;
  reg [32-1:0] _stream_matmul_16_source_7_source_ram_raddr;
  reg _stream_matmul_16_source_7_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_7_source_ram_rdata;
  reg _stream_matmul_16_source_7_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_7_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_7_source_empty_data;
  reg [1-1:0] _stream_matmul_16_parameter_8_next_parameter_data;
  reg _stream_matmul_16_source_9_idle;
  reg [33-1:0] _stream_matmul_16_source_9_source_count;
  reg [5-1:0] _stream_matmul_16_source_9_source_mode;
  reg [16-1:0] _stream_matmul_16_source_9_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_9_source_offset;
  reg [33-1:0] _stream_matmul_16_source_9_source_size;
  reg [32-1:0] _stream_matmul_16_source_9_source_stride;
  reg [32-1:0] _stream_matmul_16_source_9_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_9_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_9_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_9_source_sel;
  reg [32-1:0] _stream_matmul_16_source_9_source_ram_raddr;
  reg _stream_matmul_16_source_9_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_9_source_ram_rdata;
  reg _stream_matmul_16_source_9_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_9_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_9_source_empty_data;
  reg [1-1:0] _stream_matmul_16_parameter_10_next_parameter_data;
  reg _stream_matmul_16_source_11_idle;
  reg [33-1:0] _stream_matmul_16_source_11_source_count;
  reg [5-1:0] _stream_matmul_16_source_11_source_mode;
  reg [16-1:0] _stream_matmul_16_source_11_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_11_source_offset;
  reg [33-1:0] _stream_matmul_16_source_11_source_size;
  reg [32-1:0] _stream_matmul_16_source_11_source_stride;
  reg [32-1:0] _stream_matmul_16_source_11_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_11_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_11_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_11_source_sel;
  reg [32-1:0] _stream_matmul_16_source_11_source_ram_raddr;
  reg _stream_matmul_16_source_11_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_11_source_ram_rdata;
  reg _stream_matmul_16_source_11_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_11_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_11_source_empty_data;
  reg [1-1:0] _stream_matmul_16_parameter_12_next_parameter_data;
  reg _stream_matmul_16_source_13_idle;
  reg [33-1:0] _stream_matmul_16_source_13_source_count;
  reg [5-1:0] _stream_matmul_16_source_13_source_mode;
  reg [16-1:0] _stream_matmul_16_source_13_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_13_source_offset;
  reg [33-1:0] _stream_matmul_16_source_13_source_size;
  reg [32-1:0] _stream_matmul_16_source_13_source_stride;
  reg [32-1:0] _stream_matmul_16_source_13_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_13_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_13_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_13_source_sel;
  reg [32-1:0] _stream_matmul_16_source_13_source_ram_raddr;
  reg _stream_matmul_16_source_13_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_13_source_ram_rdata;
  reg _stream_matmul_16_source_13_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_13_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_13_source_empty_data;
  reg [1-1:0] _stream_matmul_16_parameter_14_next_parameter_data;
  reg _stream_matmul_16_source_15_idle;
  reg [33-1:0] _stream_matmul_16_source_15_source_count;
  reg [5-1:0] _stream_matmul_16_source_15_source_mode;
  reg [16-1:0] _stream_matmul_16_source_15_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_15_source_offset;
  reg [33-1:0] _stream_matmul_16_source_15_source_size;
  reg [32-1:0] _stream_matmul_16_source_15_source_stride;
  reg [32-1:0] _stream_matmul_16_source_15_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_15_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_15_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_15_source_sel;
  reg [32-1:0] _stream_matmul_16_source_15_source_ram_raddr;
  reg _stream_matmul_16_source_15_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_15_source_ram_rdata;
  reg _stream_matmul_16_source_15_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_15_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_15_source_empty_data;
  reg [1-1:0] _stream_matmul_16_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_matmul_16_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_matmul_16_parameter_18_next_parameter_data;
  reg [2-1:0] _stream_matmul_16_parameter_19_next_parameter_data;
  reg _stream_matmul_16_source_20_idle;
  reg [33-1:0] _stream_matmul_16_source_20_source_count;
  reg [5-1:0] _stream_matmul_16_source_20_source_mode;
  reg [16-1:0] _stream_matmul_16_source_20_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_20_source_offset;
  reg [33-1:0] _stream_matmul_16_source_20_source_size;
  reg [32-1:0] _stream_matmul_16_source_20_source_stride;
  reg [32-1:0] _stream_matmul_16_source_20_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_20_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_20_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_20_source_sel;
  reg [32-1:0] _stream_matmul_16_source_20_source_ram_raddr;
  reg _stream_matmul_16_source_20_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_20_source_ram_rdata;
  reg _stream_matmul_16_source_20_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_20_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_20_source_empty_data;
  reg _stream_matmul_16_source_21_idle;
  reg [33-1:0] _stream_matmul_16_source_21_source_count;
  reg [5-1:0] _stream_matmul_16_source_21_source_mode;
  reg [16-1:0] _stream_matmul_16_source_21_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_21_source_offset;
  reg [33-1:0] _stream_matmul_16_source_21_source_size;
  reg [32-1:0] _stream_matmul_16_source_21_source_stride;
  reg [32-1:0] _stream_matmul_16_source_21_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_21_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_21_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_21_source_sel;
  reg [32-1:0] _stream_matmul_16_source_21_source_ram_raddr;
  reg _stream_matmul_16_source_21_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_21_source_ram_rdata;
  reg _stream_matmul_16_source_21_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_21_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_21_source_empty_data;
  reg _stream_matmul_16_source_22_idle;
  reg [33-1:0] _stream_matmul_16_source_22_source_count;
  reg [5-1:0] _stream_matmul_16_source_22_source_mode;
  reg [16-1:0] _stream_matmul_16_source_22_source_generator_id;
  reg [32-1:0] _stream_matmul_16_source_22_source_offset;
  reg [33-1:0] _stream_matmul_16_source_22_source_size;
  reg [32-1:0] _stream_matmul_16_source_22_source_stride;
  reg [32-1:0] _stream_matmul_16_source_22_source_offset_buf;
  reg [33-1:0] _stream_matmul_16_source_22_source_size_buf;
  reg [32-1:0] _stream_matmul_16_source_22_source_stride_buf;
  reg [8-1:0] _stream_matmul_16_source_22_source_sel;
  reg [32-1:0] _stream_matmul_16_source_22_source_ram_raddr;
  reg _stream_matmul_16_source_22_source_ram_renable;
  wire [32-1:0] _stream_matmul_16_source_22_source_ram_rdata;
  reg _stream_matmul_16_source_22_source_fifo_deq;
  wire [32-1:0] _stream_matmul_16_source_22_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_16_source_22_source_empty_data;
  wire signed [64-1:0] add_tree_2_var0_data;
  wire signed [64-1:0] add_tree_2_var1_data;
  reg __add_tree_2_stream_ivalid_1;
  reg signed [64-1:0] __plusn_data_47;
  wire signed [64-1:0] add_tree_2_sum_data;
  assign add_tree_2_sum_data = __plusn_data_47;
  wire signed [64-1:0] add_tree_3_var0_data;
  wire signed [64-1:0] add_tree_3_var1_data;
  reg __add_tree_3_stream_ivalid_1;
  reg signed [64-1:0] __plusn_data_51;
  wire signed [64-1:0] add_tree_3_sum_data;
  assign add_tree_3_sum_data = __plusn_data_51;
  reg [33-1:0] _stream_matmul_16_sink_33_sink_count;
  reg [5-1:0] _stream_matmul_16_sink_33_sink_mode;
  reg [16-1:0] _stream_matmul_16_sink_33_sink_generator_id;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_offset;
  reg [33-1:0] _stream_matmul_16_sink_33_sink_size;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_stride;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_offset_buf;
  reg [33-1:0] _stream_matmul_16_sink_33_sink_size_buf;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_stride_buf;
  reg [8-1:0] _stream_matmul_16_sink_33_sink_sel;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_waddr;
  reg _stream_matmul_16_sink_33_sink_wenable;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_wdata;
  reg _stream_matmul_16_sink_33_sink_fifo_enq;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_fifo_wdata;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_immediate;
  reg [33-1:0] _stream_matmul_16_sink_34_sink_count;
  reg [5-1:0] _stream_matmul_16_sink_34_sink_mode;
  reg [16-1:0] _stream_matmul_16_sink_34_sink_generator_id;
  reg [32-1:0] _stream_matmul_16_sink_34_sink_offset;
  reg [33-1:0] _stream_matmul_16_sink_34_sink_size;
  reg [32-1:0] _stream_matmul_16_sink_34_sink_stride;
  reg [32-1:0] _stream_matmul_16_sink_34_sink_offset_buf;
  reg [33-1:0] _stream_matmul_16_sink_34_sink_size_buf;
  reg [32-1:0] _stream_matmul_16_sink_34_sink_stride_buf;
  reg [8-1:0] _stream_matmul_16_sink_34_sink_sel;
  reg [32-1:0] _stream_matmul_16_sink_34_sink_waddr;
  reg _stream_matmul_16_sink_34_sink_wenable;
  reg [1-1:0] _stream_matmul_16_sink_34_sink_wdata;
  reg _stream_matmul_16_sink_34_sink_fifo_enq;
  reg [1-1:0] _stream_matmul_16_sink_34_sink_fifo_wdata;
  reg [1-1:0] _stream_matmul_16_sink_34_sink_immediate;
  reg [32-1:0] main_fsm;
  localparam main_fsm_init = 0;
  reg [32-1:0] internal_state_counter;
  reg [32-1:0] conv2d_4_objaddr;
  reg [32-1:0] conv2d_4_arg_objaddr_0;
  reg [32-1:0] conv2d_4_arg_objaddr_1;
  reg [32-1:0] conv2d_4_arg_objaddr_2;
  reg [32-1:0] conv2d_4_arg_objaddr_3;
  reg [32-1:0] control_conv2d_4;
  localparam control_conv2d_4_init = 0;
  reg _control_conv2d_4_called;
  wire signed [32-1:0] conv2d_4_act_base_offset;
  reg signed [32-1:0] conv2d_4_act_base_offset_row;
  reg signed [32-1:0] conv2d_4_act_base_offset_bat;
  assign conv2d_4_act_base_offset = conv2d_4_act_base_offset_row + conv2d_4_act_base_offset_bat;
  reg signed [32-1:0] conv2d_4_filter_base_offset;
  reg [32-1:0] conv2d_4_next_stream_num_ops;
  wire signed [32-1:0] conv2d_4_out_base_offset;
  reg signed [32-1:0] conv2d_4_out_base_offset_val;
  reg signed [32-1:0] conv2d_4_out_base_offset_col;
  reg signed [32-1:0] conv2d_4_out_base_offset_row;
  reg signed [32-1:0] conv2d_4_out_base_offset_bat;
  reg signed [32-1:0] conv2d_4_out_base_offset_och;
  assign conv2d_4_out_base_offset = conv2d_4_out_base_offset_val + conv2d_4_out_base_offset_col + conv2d_4_out_base_offset_row + conv2d_4_out_base_offset_bat + conv2d_4_out_base_offset_och;
  reg conv2d_4_dma_flag_0;
  reg conv2d_4_dma_flag_1;
  reg conv2d_4_dma_flag_2;
  reg [32-1:0] conv2d_4_sync_comp_count;
  reg [32-1:0] conv2d_4_sync_out_count;
  reg [32-1:0] conv2d_4_write_count;
  reg [32-1:0] conv2d_4_next_out_write_size;
  reg [32-1:0] conv2d_4_col_count;
  reg [32-1:0] conv2d_4_row_count;
  reg [32-1:0] conv2d_4_bat_count;
  reg [32-1:0] conv2d_4_och_count;
  reg [2-1:0] conv2d_4_col_select;
  reg [2-1:0] conv2d_4_row_select;
  reg [32-1:0] conv2d_4_out_col_count;
  reg [32-1:0] conv2d_4_out_row_count;
  reg [32-1:0] conv2d_4_out_ram_select;
  reg [32-1:0] conv2d_4_prev_col_count;
  reg [32-1:0] conv2d_4_prev_row_count;
  reg [32-1:0] conv2d_4_prev_bat_count;
  reg [32-1:0] conv2d_4_prev_och_count;
  reg [2-1:0] conv2d_4_prev_row_select;
  reg [32-1:0] conv2d_4_stream_act_local_0;
  reg [32-1:0] conv2d_4_stream_act_local_1;
  reg [32-1:0] conv2d_4_stream_act_local_2;
  reg [32-1:0] conv2d_4_stream_act_local_3;
  reg [32-1:0] conv2d_4_stream_act_local_4;
  reg [32-1:0] conv2d_4_stream_act_local_5;
  reg [32-1:0] conv2d_4_stream_act_local_6;
  reg [32-1:0] conv2d_4_stream_act_local_7;
  reg [32-1:0] conv2d_4_stream_act_local_8;
  reg [32-1:0] conv2d_4_stream_out_local_val;
  reg [32-1:0] conv2d_4_stream_out_local_col;
  wire [32-1:0] conv2d_4_stream_out_local;
  assign conv2d_4_stream_out_local = conv2d_4_stream_out_local_val + conv2d_4_stream_out_local_col;
  reg [32-1:0] conv2d_4_act_page_comp_offset_0;
  reg [32-1:0] conv2d_4_act_page_comp_offset_1;
  reg [32-1:0] conv2d_4_act_page_comp_offset_2;
  reg [32-1:0] conv2d_4_act_page_dma_offset_0;
  reg [32-1:0] conv2d_4_act_page_dma_offset_1;
  reg [32-1:0] conv2d_4_act_page_dma_offset_2;
  reg [32-1:0] conv2d_4_filter_page_comp_offset;
  reg [32-1:0] conv2d_4_filter_page_dma_offset;
  reg conv2d_4_out_page;
  reg [32-1:0] conv2d_4_out_page_comp_offset;
  reg [32-1:0] conv2d_4_out_page_dma_offset;
  reg [32-1:0] conv2d_4_out_laddr_offset;
  reg conv2d_4_skip_read_filter;
  reg conv2d_4_skip_read_act;
  reg conv2d_4_skip_comp;
  reg conv2d_4_skip_write_out;
  wire [32-1:0] mask_addr_shifted_54;
  assign mask_addr_shifted_54 = conv2d_4_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_55;
  assign mask_addr_masked_55 = mask_addr_shifted_54 << 2;
  reg [32-1:0] _maxi_read_req_fsm;
  localparam _maxi_read_req_fsm_init = 0;
  reg [33-1:0] _maxi_read_cur_global_size;
  reg _maxi_read_cont;
  wire [8-1:0] pack_read_req_op_sel_56;
  wire [32-1:0] pack_read_req_local_addr_57;
  wire [32-1:0] pack_read_req_local_stride_58;
  wire [33-1:0] pack_read_req_local_size_59;
  wire [32-1:0] pack_read_req_local_blocksize_60;
  assign pack_read_req_op_sel_56 = _maxi_read_op_sel;
  assign pack_read_req_local_addr_57 = _maxi_read_local_addr;
  assign pack_read_req_local_stride_58 = _maxi_read_local_stride;
  assign pack_read_req_local_size_59 = _maxi_read_local_size;
  assign pack_read_req_local_blocksize_60 = _maxi_read_local_blocksize;
  wire [137-1:0] pack_read_req_packed_61;
  assign pack_read_req_packed_61 = { pack_read_req_op_sel_56, pack_read_req_local_addr_57, pack_read_req_local_stride_58, pack_read_req_local_size_59, pack_read_req_local_blocksize_60 };
  assign _maxi_read_req_fifo_wdata = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? pack_read_req_packed_61 : 'hx;
  assign _maxi_read_req_fifo_enq = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? (_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full && !_maxi_read_req_fifo_almost_full : 0;
  localparam _tmp_62 = 1;
  wire [_tmp_62-1:0] _tmp_63;
  assign _tmp_63 = !_maxi_read_req_fifo_almost_full;
  reg [_tmp_62-1:0] __tmp_63_1;
  wire [32-1:0] mask_addr_shifted_64;
  assign mask_addr_shifted_64 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_65;
  assign mask_addr_masked_65 = mask_addr_shifted_64 << 2;
  wire [32-1:0] mask_addr_shifted_66;
  assign mask_addr_shifted_66 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_67;
  assign mask_addr_masked_67 = mask_addr_shifted_66 << 2;
  wire [32-1:0] mask_addr_shifted_68;
  assign mask_addr_shifted_68 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_69;
  assign mask_addr_masked_69 = mask_addr_shifted_68 << 2;
  wire [32-1:0] mask_addr_shifted_70;
  assign mask_addr_shifted_70 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_71;
  assign mask_addr_masked_71 = mask_addr_shifted_70 << 2;
  wire [32-1:0] mask_addr_shifted_72;
  assign mask_addr_shifted_72 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_73;
  assign mask_addr_masked_73 = mask_addr_shifted_72 << 2;
  wire [32-1:0] mask_addr_shifted_74;
  assign mask_addr_shifted_74 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_75;
  assign mask_addr_masked_75 = mask_addr_shifted_74 << 2;
  reg _maxi_raddr_cond_0_1;
  reg [32-1:0] _maxi_read_data_fsm;
  localparam _maxi_read_data_fsm_init = 0;
  reg [32-1:0] write_burst_fsm_0;
  localparam write_burst_fsm_0_init = 0;
  reg [7-1:0] write_burst_addr_76;
  reg [7-1:0] write_burst_stride_77;
  reg [33-1:0] write_burst_length_78;
  reg write_burst_done_79;
  assign ram_w32_l128_id18_1_addr = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_76 : 'hx;
  assign ram_w32_l128_id18_1_wdata = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id18_1_wenable = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l128_id18_1_enable = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_80;
  assign mask_addr_shifted_80 = conv2d_4_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_81;
  assign mask_addr_masked_81 = mask_addr_shifted_80 << 2;
  reg [32-1:0] write_burst_fsm_1;
  localparam write_burst_fsm_1_init = 0;
  reg [7-1:0] write_burst_addr_82;
  reg [7-1:0] write_burst_stride_83;
  reg [33-1:0] write_burst_length_84;
  reg write_burst_done_85;
  assign ram_w32_l128_id19_1_addr = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_82 : 'hx;
  assign ram_w32_l128_id19_1_wdata = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id19_1_wenable = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l128_id19_1_enable = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_86;
  assign mask_addr_shifted_86 = conv2d_4_arg_objaddr_1 + conv2d_4_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_87;
  assign mask_addr_masked_87 = mask_addr_shifted_86 << 2;
  wire write_burst_block_ram_wvalid_88;
  wire write_burst_block_ram_wquit_89;
  reg [32-1:0] write_burst_fsm_2;
  localparam write_burst_fsm_2_init = 0;
  reg [7-1:0] write_burst_addr_90;
  reg [7-1:0] write_burst_stride_91;
  reg [33-1:0] write_burst_length_92;
  reg write_burst_done_93;
  assign ram_w32_l128_id0_1_wdata = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id0_1_wenable = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_94;
  wire write_burst_block_ram_wquit_95;
  reg [32-1:0] write_burst_fsm_3;
  localparam write_burst_fsm_3_init = 0;
  reg [7-1:0] write_burst_addr_96;
  reg [7-1:0] write_burst_stride_97;
  reg [33-1:0] write_burst_length_98;
  reg write_burst_done_99;
  assign ram_w32_l128_id1_1_addr = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? write_burst_addr_96 : 'hx;
  assign ram_w32_l128_id1_1_wdata = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id1_1_wenable = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? 1'd1 : 0;
  assign ram_w32_l128_id1_1_enable = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_100;
  wire write_burst_block_ram_wquit_101;
  reg [32-1:0] write_burst_fsm_4;
  localparam write_burst_fsm_4_init = 0;
  reg [7-1:0] write_burst_addr_102;
  reg [7-1:0] write_burst_stride_103;
  reg [33-1:0] write_burst_length_104;
  reg write_burst_done_105;
  assign ram_w32_l128_id2_1_addr = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? write_burst_addr_102 : 'hx;
  assign ram_w32_l128_id2_1_wdata = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id2_1_wenable = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? 1'd1 : 0;
  assign ram_w32_l128_id2_1_enable = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_106;
  wire write_burst_block_ram_wquit_107;
  reg [32-1:0] write_burst_fsm_5;
  localparam write_burst_fsm_5_init = 0;
  reg [7-1:0] write_burst_addr_108;
  reg [7-1:0] write_burst_stride_109;
  reg [33-1:0] write_burst_length_110;
  reg write_burst_done_111;
  assign ram_w32_l128_id3_1_addr = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? write_burst_addr_108 : 'hx;
  assign ram_w32_l128_id3_1_wdata = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id3_1_wenable = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? 1'd1 : 0;
  assign ram_w32_l128_id3_1_enable = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_112;
  wire write_burst_block_ram_wquit_113;
  reg [32-1:0] write_burst_fsm_6;
  localparam write_burst_fsm_6_init = 0;
  reg [7-1:0] write_burst_addr_114;
  reg [7-1:0] write_burst_stride_115;
  reg [33-1:0] write_burst_length_116;
  reg write_burst_done_117;
  assign ram_w32_l128_id4_1_addr = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? write_burst_addr_114 : 'hx;
  assign ram_w32_l128_id4_1_wdata = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id4_1_wenable = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? 1'd1 : 0;
  assign ram_w32_l128_id4_1_enable = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_118;
  wire write_burst_block_ram_wquit_119;
  reg [32-1:0] write_burst_fsm_7;
  localparam write_burst_fsm_7_init = 0;
  reg [7-1:0] write_burst_addr_120;
  reg [7-1:0] write_burst_stride_121;
  reg [33-1:0] write_burst_length_122;
  reg write_burst_done_123;
  assign ram_w32_l128_id5_1_addr = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? write_burst_addr_120 : 'hx;
  assign ram_w32_l128_id5_1_wdata = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id5_1_wenable = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  assign ram_w32_l128_id5_1_enable = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_124;
  wire write_burst_block_ram_wquit_125;
  reg [32-1:0] write_burst_fsm_8;
  localparam write_burst_fsm_8_init = 0;
  reg [7-1:0] write_burst_addr_126;
  reg [7-1:0] write_burst_stride_127;
  reg [33-1:0] write_burst_length_128;
  reg write_burst_done_129;
  assign ram_w32_l128_id6_1_addr = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? write_burst_addr_126 : 'hx;
  assign ram_w32_l128_id6_1_wdata = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id6_1_wenable = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? 1'd1 : 0;
  assign ram_w32_l128_id6_1_enable = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_130;
  wire write_burst_block_ram_wquit_131;
  reg [32-1:0] write_burst_fsm_9;
  localparam write_burst_fsm_9_init = 0;
  reg [7-1:0] write_burst_addr_132;
  reg [7-1:0] write_burst_stride_133;
  reg [33-1:0] write_burst_length_134;
  reg write_burst_done_135;
  assign ram_w32_l128_id7_1_addr = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? write_burst_addr_132 : 'hx;
  assign ram_w32_l128_id7_1_wdata = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id7_1_wenable = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? 1'd1 : 0;
  assign ram_w32_l128_id7_1_enable = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_136;
  wire write_burst_block_ram_wquit_137;
  reg [32-1:0] write_burst_fsm_10;
  localparam write_burst_fsm_10_init = 0;
  reg [7-1:0] write_burst_addr_138;
  reg [7-1:0] write_burst_stride_139;
  reg [33-1:0] write_burst_length_140;
  reg write_burst_done_141;
  assign ram_w32_l128_id8_1_addr = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? write_burst_addr_138 : 'hx;
  assign ram_w32_l128_id8_1_wdata = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id8_1_wenable = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? 1'd1 : 0;
  assign ram_w32_l128_id8_1_enable = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_142;
  wire write_burst_block_ram_wquit_143;
  reg [32-1:0] write_burst_fsm_11;
  localparam write_burst_fsm_11_init = 0;
  reg [7-1:0] write_burst_addr_144;
  reg [7-1:0] write_burst_stride_145;
  reg [33-1:0] write_burst_length_146;
  reg write_burst_done_147;
  assign ram_w32_l128_id9_1_addr = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_142)? write_burst_addr_144 : 'hx;
  assign ram_w32_l128_id9_1_wdata = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_142)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id9_1_wenable = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_142)? 1'd1 : 0;
  assign ram_w32_l128_id9_1_enable = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_142)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_148;
  wire write_burst_block_ram_wquit_149;
  reg [32-1:0] write_burst_fsm_12;
  localparam write_burst_fsm_12_init = 0;
  reg [7-1:0] write_burst_addr_150;
  reg [7-1:0] write_burst_stride_151;
  reg [33-1:0] write_burst_length_152;
  reg write_burst_done_153;
  assign ram_w32_l128_id10_1_addr = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? write_burst_addr_150 : 'hx;
  assign ram_w32_l128_id10_1_wdata = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id10_1_wenable = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  assign ram_w32_l128_id10_1_enable = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_154;
  wire write_burst_block_ram_wquit_155;
  reg [32-1:0] write_burst_fsm_13;
  localparam write_burst_fsm_13_init = 0;
  reg [7-1:0] write_burst_addr_156;
  reg [7-1:0] write_burst_stride_157;
  reg [33-1:0] write_burst_length_158;
  reg write_burst_done_159;
  assign ram_w32_l128_id11_1_addr = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? write_burst_addr_156 : 'hx;
  assign ram_w32_l128_id11_1_wdata = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id11_1_wenable = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? 1'd1 : 0;
  assign ram_w32_l128_id11_1_enable = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_160;
  wire write_burst_block_ram_wquit_161;
  reg [32-1:0] write_burst_fsm_14;
  localparam write_burst_fsm_14_init = 0;
  reg [7-1:0] write_burst_addr_162;
  reg [7-1:0] write_burst_stride_163;
  reg [33-1:0] write_burst_length_164;
  reg write_burst_done_165;
  assign ram_w32_l128_id12_1_addr = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? write_burst_addr_162 : 'hx;
  assign ram_w32_l128_id12_1_wdata = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id12_1_wenable = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? 1'd1 : 0;
  assign ram_w32_l128_id12_1_enable = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_166;
  wire write_burst_block_ram_wquit_167;
  reg [32-1:0] write_burst_fsm_15;
  localparam write_burst_fsm_15_init = 0;
  reg [7-1:0] write_burst_addr_168;
  reg [7-1:0] write_burst_stride_169;
  reg [33-1:0] write_burst_length_170;
  reg write_burst_done_171;
  assign ram_w32_l128_id13_1_addr = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_166)? write_burst_addr_168 : 'hx;
  assign ram_w32_l128_id13_1_wdata = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_166)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id13_1_wenable = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_166)? 1'd1 : 0;
  assign ram_w32_l128_id13_1_enable = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_166)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_172;
  wire write_burst_block_ram_wquit_173;
  reg [32-1:0] write_burst_fsm_16;
  localparam write_burst_fsm_16_init = 0;
  reg [7-1:0] write_burst_addr_174;
  reg [7-1:0] write_burst_stride_175;
  reg [33-1:0] write_burst_length_176;
  reg write_burst_done_177;
  assign ram_w32_l128_id14_1_addr = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? write_burst_addr_174 : 'hx;
  assign ram_w32_l128_id14_1_wdata = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id14_1_wenable = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? 1'd1 : 0;
  assign ram_w32_l128_id14_1_enable = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_178;
  wire write_burst_block_ram_wquit_179;
  reg [32-1:0] write_burst_fsm_17;
  localparam write_burst_fsm_17_init = 0;
  reg [7-1:0] write_burst_addr_180;
  reg [7-1:0] write_burst_stride_181;
  reg [33-1:0] write_burst_length_182;
  reg write_burst_done_183;
  assign ram_w32_l128_id15_1_addr = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? write_burst_addr_180 : 'hx;
  assign ram_w32_l128_id15_1_wdata = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id15_1_wenable = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  assign ram_w32_l128_id15_1_enable = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_184;
  wire write_burst_block_ram_wquit_185;
  reg [32-1:0] write_burst_fsm_18;
  localparam write_burst_fsm_18_init = 0;
  reg [7-1:0] write_burst_addr_186;
  reg [7-1:0] write_burst_stride_187;
  reg [33-1:0] write_burst_length_188;
  reg write_burst_done_189;
  assign ram_w32_l128_id16_1_addr = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? write_burst_addr_186 : 'hx;
  assign ram_w32_l128_id16_1_wdata = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id16_1_wenable = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? 1'd1 : 0;
  assign ram_w32_l128_id16_1_enable = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_190;
  wire write_burst_block_ram_wquit_191;
  reg [32-1:0] write_burst_fsm_19;
  localparam write_burst_fsm_19_init = 0;
  reg [7-1:0] write_burst_addr_192;
  reg [7-1:0] write_burst_stride_193;
  reg [33-1:0] write_burst_length_194;
  reg write_burst_done_195;
  assign ram_w32_l128_id17_1_addr = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_190)? write_burst_addr_192 : 'hx;
  assign ram_w32_l128_id17_1_wdata = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_190)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l128_id17_1_wenable = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_190)? 1'd1 : 0;
  assign ram_w32_l128_id17_1_enable = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_190)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_20;
  localparam write_burst_block_fsm_20_init = 0;
  reg [33-1:0] write_burst_block_length_196;
  reg [32-1:0] write_burst_block_blocksize_197;
  reg write_burst_block_done_198;
  reg [32-1:0] write_burst_block_count_199;
  assign write_burst_block_ram_wvalid_88 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 1);
  assign write_burst_block_ram_wquit_89 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_94 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 2);
  assign write_burst_block_ram_wquit_95 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_100 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 3);
  assign write_burst_block_ram_wquit_101 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_106 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 4);
  assign write_burst_block_ram_wquit_107 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_112 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 5);
  assign write_burst_block_ram_wquit_113 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_118 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 6);
  assign write_burst_block_ram_wquit_119 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_124 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 7);
  assign write_burst_block_ram_wquit_125 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_130 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 8);
  assign write_burst_block_ram_wquit_131 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_136 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 9);
  assign write_burst_block_ram_wquit_137 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_142 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 10);
  assign write_burst_block_ram_wquit_143 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_148 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 11);
  assign write_burst_block_ram_wquit_149 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_154 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 12);
  assign write_burst_block_ram_wquit_155 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_160 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 13);
  assign write_burst_block_ram_wquit_161 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_166 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 14);
  assign write_burst_block_ram_wquit_167 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_172 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 15);
  assign write_burst_block_ram_wquit_173 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_178 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 16);
  assign write_burst_block_ram_wquit_179 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_184 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 17);
  assign write_burst_block_ram_wquit_185 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  assign write_burst_block_ram_wvalid_190 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_20 == 18);
  assign write_burst_block_ram_wquit_191 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1);
  wire [32-1:0] conv2d_4_mux_act_gaddr_0;
  assign conv2d_4_mux_act_gaddr_0 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 1'd0;
  wire [32-1:0] conv2d_4_mux_act_gaddr_1;
  assign conv2d_4_mux_act_gaddr_1 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 1'd0;
  wire [32-1:0] conv2d_4_mux_act_gaddr_2;
  assign conv2d_4_mux_act_gaddr_2 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 1'd0;
  wire conv2d_4_dma_pad_mask_0;
  assign conv2d_4_dma_pad_mask_0 = (conv2d_4_row_count + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_dma_pad_mask_1;
  assign conv2d_4_dma_pad_mask_1 = (conv2d_4_row_count + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_dma_pad_mask_2;
  assign conv2d_4_dma_pad_mask_2 = (conv2d_4_row_count + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_mux_dma_pad_mask_0;
  assign conv2d_4_mux_dma_pad_mask_0 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_0 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_2 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_1 : 1'd0;
  wire conv2d_4_mux_dma_pad_mask_1;
  assign conv2d_4_mux_dma_pad_mask_1 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_1 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_0 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_2 : 1'd0;
  wire conv2d_4_mux_dma_pad_mask_2;
  assign conv2d_4_mux_dma_pad_mask_2 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_2 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_1 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_0 : 1'd0;
  wire conv2d_4_mux_dma_flag_0;
  assign conv2d_4_mux_dma_flag_0 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_0 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_2 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_1 : 1'd0;
  wire conv2d_4_mux_dma_flag_1;
  assign conv2d_4_mux_dma_flag_1 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_1 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_0 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_2 : 1'd0;
  wire conv2d_4_mux_dma_flag_2;
  assign conv2d_4_mux_dma_flag_2 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_2 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_1 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_0 : 1'd0;
  wire [32-1:0] mask_addr_shifted_200;
  assign mask_addr_shifted_200 = conv2d_4_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_201;
  assign mask_addr_masked_201 = mask_addr_shifted_200 << 2;
  wire write_burst_block_ram_wvalid_202;
  wire write_burst_block_ram_wquit_203;
  reg [32-1:0] write_burst_fsm_21;
  localparam write_burst_fsm_21_init = 0;
  reg [9-1:0] write_burst_addr_204;
  reg [9-1:0] write_burst_stride_205;
  reg [33-1:0] write_burst_length_206;
  reg write_burst_done_207;
  assign ram_w32_l512_id0_1_addr = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? write_burst_addr_204 : 'hx;
  assign ram_w32_l512_id0_1_wdata = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id0_1_wenable = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? 1'd1 : 0;
  assign ram_w32_l512_id0_1_enable = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_208;
  wire write_burst_block_ram_wquit_209;
  reg [32-1:0] write_burst_fsm_22;
  localparam write_burst_fsm_22_init = 0;
  reg [9-1:0] write_burst_addr_210;
  reg [9-1:0] write_burst_stride_211;
  reg [33-1:0] write_burst_length_212;
  reg write_burst_done_213;
  assign ram_w32_l512_id1_1_addr = ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? write_burst_addr_210 : 'hx;
  assign ram_w32_l512_id1_1_wdata = ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id1_1_wenable = ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? 1'd1 : 0;
  assign ram_w32_l512_id1_1_enable = ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_214;
  wire write_burst_block_ram_wquit_215;
  reg [32-1:0] write_burst_fsm_23;
  localparam write_burst_fsm_23_init = 0;
  reg [9-1:0] write_burst_addr_216;
  reg [9-1:0] write_burst_stride_217;
  reg [33-1:0] write_burst_length_218;
  reg write_burst_done_219;
  assign ram_w32_l512_id2_1_addr = ((write_burst_fsm_23 == 1) && write_burst_block_ram_wvalid_214)? write_burst_addr_216 : 'hx;
  assign ram_w32_l512_id2_1_wdata = ((write_burst_fsm_23 == 1) && write_burst_block_ram_wvalid_214)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id2_1_wenable = ((write_burst_fsm_23 == 1) && write_burst_block_ram_wvalid_214)? 1'd1 : 0;
  assign ram_w32_l512_id2_1_enable = ((write_burst_fsm_23 == 1) && write_burst_block_ram_wvalid_214)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_24;
  localparam write_burst_block_fsm_24_init = 0;
  reg [33-1:0] write_burst_block_length_220;
  reg [32-1:0] write_burst_block_blocksize_221;
  reg write_burst_block_done_222;
  reg [32-1:0] write_burst_block_count_223;
  assign write_burst_block_ram_wvalid_202 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_24 == 1);
  assign write_burst_block_ram_wquit_203 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1);
  assign write_burst_block_ram_wvalid_208 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_24 == 2);
  assign write_burst_block_ram_wquit_209 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1);
  assign write_burst_block_ram_wvalid_214 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_24 == 3);
  assign write_burst_block_ram_wquit_215 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1);
  wire [32-1:0] mask_addr_shifted_224;
  assign mask_addr_shifted_224 = conv2d_4_mux_act_gaddr_1 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_225;
  assign mask_addr_masked_225 = mask_addr_shifted_224 << 2;
  wire write_burst_block_ram_wvalid_226;
  wire write_burst_block_ram_wquit_227;
  reg [32-1:0] write_burst_fsm_25;
  localparam write_burst_fsm_25_init = 0;
  reg [9-1:0] write_burst_addr_228;
  reg [9-1:0] write_burst_stride_229;
  reg [33-1:0] write_burst_length_230;
  reg write_burst_done_231;
  assign ram_w32_l512_id3_1_addr = ((write_burst_fsm_25 == 1) && write_burst_block_ram_wvalid_226)? write_burst_addr_228 : 'hx;
  assign ram_w32_l512_id3_1_wdata = ((write_burst_fsm_25 == 1) && write_burst_block_ram_wvalid_226)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id3_1_wenable = ((write_burst_fsm_25 == 1) && write_burst_block_ram_wvalid_226)? 1'd1 : 0;
  assign ram_w32_l512_id3_1_enable = ((write_burst_fsm_25 == 1) && write_burst_block_ram_wvalid_226)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_232;
  wire write_burst_block_ram_wquit_233;
  reg [32-1:0] write_burst_fsm_26;
  localparam write_burst_fsm_26_init = 0;
  reg [9-1:0] write_burst_addr_234;
  reg [9-1:0] write_burst_stride_235;
  reg [33-1:0] write_burst_length_236;
  reg write_burst_done_237;
  assign ram_w32_l512_id4_1_addr = ((write_burst_fsm_26 == 1) && write_burst_block_ram_wvalid_232)? write_burst_addr_234 : 'hx;
  assign ram_w32_l512_id4_1_wdata = ((write_burst_fsm_26 == 1) && write_burst_block_ram_wvalid_232)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id4_1_wenable = ((write_burst_fsm_26 == 1) && write_burst_block_ram_wvalid_232)? 1'd1 : 0;
  assign ram_w32_l512_id4_1_enable = ((write_burst_fsm_26 == 1) && write_burst_block_ram_wvalid_232)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_238;
  wire write_burst_block_ram_wquit_239;
  reg [32-1:0] write_burst_fsm_27;
  localparam write_burst_fsm_27_init = 0;
  reg [9-1:0] write_burst_addr_240;
  reg [9-1:0] write_burst_stride_241;
  reg [33-1:0] write_burst_length_242;
  reg write_burst_done_243;
  assign ram_w32_l512_id5_1_addr = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_238)? write_burst_addr_240 : 'hx;
  assign ram_w32_l512_id5_1_wdata = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_238)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id5_1_wenable = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_238)? 1'd1 : 0;
  assign ram_w32_l512_id5_1_enable = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_238)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_28;
  localparam write_burst_block_fsm_28_init = 0;
  reg [33-1:0] write_burst_block_length_244;
  reg [32-1:0] write_burst_block_blocksize_245;
  reg write_burst_block_done_246;
  reg [32-1:0] write_burst_block_count_247;
  assign write_burst_block_ram_wvalid_226 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_28 == 1);
  assign write_burst_block_ram_wquit_227 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1);
  assign write_burst_block_ram_wvalid_232 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_28 == 2);
  assign write_burst_block_ram_wquit_233 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1);
  assign write_burst_block_ram_wvalid_238 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_28 == 3);
  assign write_burst_block_ram_wquit_239 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1);
  wire [32-1:0] mask_addr_shifted_248;
  assign mask_addr_shifted_248 = conv2d_4_mux_act_gaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_249;
  assign mask_addr_masked_249 = mask_addr_shifted_248 << 2;
  wire write_burst_block_ram_wvalid_250;
  wire write_burst_block_ram_wquit_251;
  reg [32-1:0] write_burst_fsm_29;
  localparam write_burst_fsm_29_init = 0;
  reg [9-1:0] write_burst_addr_252;
  reg [9-1:0] write_burst_stride_253;
  reg [33-1:0] write_burst_length_254;
  reg write_burst_done_255;
  assign ram_w32_l512_id6_1_addr = ((write_burst_fsm_29 == 1) && write_burst_block_ram_wvalid_250)? write_burst_addr_252 : 'hx;
  assign ram_w32_l512_id6_1_wdata = ((write_burst_fsm_29 == 1) && write_burst_block_ram_wvalid_250)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id6_1_wenable = ((write_burst_fsm_29 == 1) && write_burst_block_ram_wvalid_250)? 1'd1 : 0;
  assign ram_w32_l512_id6_1_enable = ((write_burst_fsm_29 == 1) && write_burst_block_ram_wvalid_250)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_256;
  wire write_burst_block_ram_wquit_257;
  reg [32-1:0] write_burst_fsm_30;
  localparam write_burst_fsm_30_init = 0;
  reg [9-1:0] write_burst_addr_258;
  reg [9-1:0] write_burst_stride_259;
  reg [33-1:0] write_burst_length_260;
  reg write_burst_done_261;
  assign ram_w32_l512_id7_1_addr = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_256)? write_burst_addr_258 : 'hx;
  assign ram_w32_l512_id7_1_wdata = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_256)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id7_1_wenable = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_256)? 1'd1 : 0;
  assign ram_w32_l512_id7_1_enable = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_256)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_262;
  wire write_burst_block_ram_wquit_263;
  reg [32-1:0] write_burst_fsm_31;
  localparam write_burst_fsm_31_init = 0;
  reg [9-1:0] write_burst_addr_264;
  reg [9-1:0] write_burst_stride_265;
  reg [33-1:0] write_burst_length_266;
  reg write_burst_done_267;
  assign ram_w32_l512_id8_1_addr = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_262)? write_burst_addr_264 : 'hx;
  assign ram_w32_l512_id8_1_wdata = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_262)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l512_id8_1_wenable = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  assign ram_w32_l512_id8_1_enable = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_32;
  localparam write_burst_block_fsm_32_init = 0;
  reg [33-1:0] write_burst_block_length_268;
  reg [32-1:0] write_burst_block_blocksize_269;
  reg write_burst_block_done_270;
  reg [32-1:0] write_burst_block_count_271;
  assign write_burst_block_ram_wvalid_250 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_32 == 1);
  assign write_burst_block_ram_wquit_251 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1);
  assign write_burst_block_ram_wvalid_256 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_32 == 2);
  assign write_burst_block_ram_wquit_257 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1);
  assign write_burst_block_ram_wvalid_262 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_32 == 3);
  assign write_burst_block_ram_wquit_263 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1);
  reg [32-1:0] conv2d_4_comp_fsm;
  localparam conv2d_4_comp_fsm_init = 0;
  reg [32-1:0] conv2d_4_filter_page_comp_offset_buf;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_0;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_1;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_2;
  reg [32-1:0] conv2d_4_out_page_comp_offset_buf;
  reg [32-1:0] conv2d_4_row_count_buf;
  reg [2-1:0] conv2d_4_row_select_buf;
  reg [32-1:0] conv2d_4_och_count_buf;
  wire conv2d_4_stream_pad_mask_0_0;
  assign conv2d_4_stream_pad_mask_0_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_0_1;
  assign conv2d_4_stream_pad_mask_0_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_0_2;
  assign conv2d_4_stream_pad_mask_0_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_0;
  assign conv2d_4_stream_pad_mask_1_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_1;
  assign conv2d_4_stream_pad_mask_1_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_2;
  assign conv2d_4_stream_pad_mask_1_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_0;
  assign conv2d_4_stream_pad_mask_2_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_1;
  assign conv2d_4_stream_pad_mask_2_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_2;
  assign conv2d_4_stream_pad_mask_2_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  reg [9-1:0] conv2d_4_stream_pad_masks;
  wire [6-1:0] stream_conv2d_4_parameter_0_data;
  wire [2-1:0] stream_conv2d_4_parameter_1_data;
  wire [2-1:0] stream_conv2d_4_parameter_2_data;
  wire [9-1:0] stream_conv2d_4_parameter_3_data;
  wire [2-1:0] stream_conv2d_4_parameter_4_data;
  wire [1-1:0] stream_conv2d_4__reduce_reset_data;
  wire [1-1:0] stream_conv2d_4_parameter_6_data;
  wire [32-1:0] stream_conv2d_4_source_7_data;
  wire [1-1:0] stream_conv2d_4_parameter_8_data;
  wire [32-1:0] stream_conv2d_4_source_9_data;
  wire [1-1:0] stream_conv2d_4_parameter_10_data;
  wire [32-1:0] stream_conv2d_4_source_11_data;
  wire [1-1:0] stream_conv2d_4_parameter_12_data;
  wire [32-1:0] stream_conv2d_4_source_13_data;
  wire [1-1:0] stream_conv2d_4_parameter_14_data;
  wire [32-1:0] stream_conv2d_4_source_15_data;
  wire [1-1:0] stream_conv2d_4_parameter_16_data;
  wire [1-1:0] stream_conv2d_4_parameter_17_data;
  wire [5-1:0] stream_conv2d_4_parameter_18_data;
  wire [1-1:0] stream_conv2d_4_parameter_19_data;
  wire [32-1:0] stream_conv2d_4_source_20_data;
  wire [32-1:0] stream_conv2d_4_source_21_data;
  wire [32-1:0] stream_conv2d_4_source_22_data;
  wire [32-1:0] stream_conv2d_4_source_23_data;
  wire [32-1:0] stream_conv2d_4_source_24_data;
  wire [32-1:0] stream_conv2d_4_source_25_data;
  wire [32-1:0] stream_conv2d_4_source_26_data;
  wire [32-1:0] stream_conv2d_4_source_27_data;
  wire [32-1:0] stream_conv2d_4_source_28_data;
  wire [32-1:0] stream_conv2d_4_source_29_data;
  wire [32-1:0] stream_conv2d_4_source_30_data;
  wire [32-1:0] stream_conv2d_4_source_31_data;
  wire [32-1:0] stream_conv2d_4_source_32_data;
  wire [32-1:0] stream_conv2d_4_source_33_data;
  wire [32-1:0] stream_conv2d_4_source_34_data;
  wire [32-1:0] stream_conv2d_4_source_35_data;
  wire [32-1:0] stream_conv2d_4_source_36_data;
  wire [32-1:0] stream_conv2d_4_source_37_data;
  wire [32-1:0] stream_conv2d_4_source_38_data;
  wire [32-1:0] stream_conv2d_4_source_39_data;
  wire [32-1:0] stream_conv2d_4_source_40_data;
  wire [32-1:0] stream_conv2d_4_source_41_data;
  wire [32-1:0] stream_conv2d_4_source_42_data;
  wire [32-1:0] stream_conv2d_4_source_43_data;
  wire [32-1:0] stream_conv2d_4_source_44_data;
  wire [32-1:0] stream_conv2d_4_source_45_data;
  wire [32-1:0] stream_conv2d_4_source_46_data;
  reg __stream_conv2d_4_stream_ivalid_1;
  reg __stream_conv2d_4_stream_ivalid_2;
  reg __stream_conv2d_4_stream_ivalid_3;
  reg __stream_conv2d_4_stream_ivalid_4;
  reg __stream_conv2d_4_stream_ivalid_5;
  reg __stream_conv2d_4_stream_ivalid_6;
  reg __stream_conv2d_4_stream_ivalid_7;
  reg __stream_conv2d_4_stream_ivalid_8;
  reg __stream_conv2d_4_stream_ivalid_9;
  reg __stream_conv2d_4_stream_ivalid_10;
  reg __stream_conv2d_4_stream_ivalid_11;
  reg __stream_conv2d_4_stream_ivalid_12;
  reg __stream_conv2d_4_stream_ivalid_13;
  reg __stream_conv2d_4_stream_ivalid_14;
  reg __stream_conv2d_4_stream_ivalid_15;
  reg __stream_conv2d_4_stream_ivalid_16;
  reg __stream_conv2d_4_stream_ivalid_17;
  reg __stream_conv2d_4_stream_ivalid_18;
  reg __stream_conv2d_4_stream_ivalid_19;
  reg __stream_conv2d_4_stream_ivalid_20;
  reg __stream_conv2d_4_stream_ivalid_21;
  reg __stream_conv2d_4_stream_ivalid_22;
  reg __stream_conv2d_4_stream_ivalid_23;
  reg __stream_conv2d_4_stream_ivalid_24;
  reg __stream_conv2d_4_stream_ivalid_25;
  reg __stream_conv2d_4_stream_ivalid_26;
  reg __stream_conv2d_4_stream_ivalid_27;
  reg __stream_conv2d_4_stream_ivalid_28;
  reg __stream_conv2d_4_stream_ivalid_29;
  reg __stream_conv2d_4_stream_ivalid_30;
  reg __stream_conv2d_4_stream_ivalid_31;
  reg __stream_conv2d_4_stream_ivalid_32;
  reg __stream_conv2d_4_stream_ivalid_33;
  reg __stream_conv2d_4_stream_ivalid_34;
  reg [32-1:0] _counter_data_952;
  reg [32-1:0] _counter_count_952;
  wire _counter_reset_cond_952;
  assign _counter_reset_cond_952 = stream_conv2d_4__reduce_reset_data;
  wire [32-1:0] _counter_current_count_952;
  assign _counter_current_count_952 = (_counter_reset_cond_952)? 1'sd0 : _counter_count_952;
  wire [1-1:0] _pointer_data_955;
  assign _pointer_data_955 = stream_conv2d_4_parameter_4_data[1'sd0];
  reg [6-1:0] _minus_data_957;
  wire [1-1:0] _pointer_data_961;
  assign _pointer_data_961 = stream_conv2d_4_parameter_4_data[2'sd1];
  reg [6-1:0] _minus_data_963;
  wire [16-1:0] _slice_data_971;
  assign _slice_data_971 = stream_conv2d_4_source_7_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_972;
  assign _reinterpretcast_src_972 = _slice_data_971;
  wire signed [16-1:0] _reinterpretcast_data_972;
  assign _reinterpretcast_data_972 = _reinterpretcast_src_972;
  wire [16-1:0] _slice_data_975;
  assign _slice_data_975 = stream_conv2d_4_source_7_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_976;
  assign _reinterpretcast_src_976 = _slice_data_975;
  wire signed [16-1:0] _reinterpretcast_data_976;
  assign _reinterpretcast_data_976 = _reinterpretcast_src_976;
  wire signed [16-1:0] _cond_data_977;
  assign _cond_data_977 = (stream_conv2d_4_parameter_6_data)? _reinterpretcast_data_972 : _reinterpretcast_data_972;
  wire signed [16-1:0] _cond_data_978;
  assign _cond_data_978 = (stream_conv2d_4_parameter_6_data)? _reinterpretcast_data_972 : _reinterpretcast_data_976;
  wire [16-1:0] _slice_data_983;
  assign _slice_data_983 = stream_conv2d_4_source_9_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_984;
  assign _reinterpretcast_src_984 = _slice_data_983;
  wire signed [16-1:0] _reinterpretcast_data_984;
  assign _reinterpretcast_data_984 = _reinterpretcast_src_984;
  wire [16-1:0] _slice_data_987;
  assign _slice_data_987 = stream_conv2d_4_source_9_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_988;
  assign _reinterpretcast_src_988 = _slice_data_987;
  wire signed [16-1:0] _reinterpretcast_data_988;
  assign _reinterpretcast_data_988 = _reinterpretcast_src_988;
  wire signed [16-1:0] _cond_data_989;
  assign _cond_data_989 = (stream_conv2d_4_parameter_8_data)? _reinterpretcast_data_984 : _reinterpretcast_data_984;
  wire signed [16-1:0] _cond_data_990;
  assign _cond_data_990 = (stream_conv2d_4_parameter_8_data)? _reinterpretcast_data_984 : _reinterpretcast_data_988;
  wire [16-1:0] _slice_data_995;
  assign _slice_data_995 = stream_conv2d_4_source_11_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_996;
  assign _reinterpretcast_src_996 = _slice_data_995;
  wire [16-1:0] _reinterpretcast_data_996;
  assign _reinterpretcast_data_996 = _reinterpretcast_src_996;
  wire [16-1:0] _slice_data_999;
  assign _slice_data_999 = stream_conv2d_4_source_11_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1000;
  assign _reinterpretcast_src_1000 = _slice_data_999;
  wire [16-1:0] _reinterpretcast_data_1000;
  assign _reinterpretcast_data_1000 = _reinterpretcast_src_1000;
  wire [16-1:0] _cond_data_1001;
  assign _cond_data_1001 = (stream_conv2d_4_parameter_10_data)? _reinterpretcast_data_996 : _reinterpretcast_data_996;
  wire [16-1:0] _cond_data_1002;
  assign _cond_data_1002 = (stream_conv2d_4_parameter_10_data)? _reinterpretcast_data_996 : _reinterpretcast_data_1000;
  wire [16-1:0] _slice_data_1007;
  assign _slice_data_1007 = stream_conv2d_4_source_13_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1008;
  assign _reinterpretcast_src_1008 = _slice_data_1007;
  wire [16-1:0] _reinterpretcast_data_1008;
  assign _reinterpretcast_data_1008 = _reinterpretcast_src_1008;
  wire [16-1:0] _slice_data_1011;
  assign _slice_data_1011 = stream_conv2d_4_source_13_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1012;
  assign _reinterpretcast_src_1012 = _slice_data_1011;
  wire [16-1:0] _reinterpretcast_data_1012;
  assign _reinterpretcast_data_1012 = _reinterpretcast_src_1012;
  wire [16-1:0] _cond_data_1013;
  assign _cond_data_1013 = (stream_conv2d_4_parameter_12_data)? _reinterpretcast_data_1008 : _reinterpretcast_data_1008;
  wire [16-1:0] _cond_data_1014;
  assign _cond_data_1014 = (stream_conv2d_4_parameter_12_data)? _reinterpretcast_data_1008 : _reinterpretcast_data_1012;
  wire [16-1:0] _slice_data_1019;
  assign _slice_data_1019 = stream_conv2d_4_source_15_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1020;
  assign _reinterpretcast_src_1020 = _slice_data_1019;
  wire [16-1:0] _reinterpretcast_data_1020;
  assign _reinterpretcast_data_1020 = _reinterpretcast_src_1020;
  wire [16-1:0] _slice_data_1023;
  assign _slice_data_1023 = stream_conv2d_4_source_15_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1024;
  assign _reinterpretcast_src_1024 = _slice_data_1023;
  wire [16-1:0] _reinterpretcast_data_1024;
  assign _reinterpretcast_data_1024 = _reinterpretcast_src_1024;
  wire [16-1:0] _cond_data_1025;
  assign _cond_data_1025 = (stream_conv2d_4_parameter_14_data)? _reinterpretcast_data_1020 : _reinterpretcast_data_1020;
  wire [16-1:0] _cond_data_1026;
  assign _cond_data_1026 = (stream_conv2d_4_parameter_14_data)? _reinterpretcast_data_1020 : _reinterpretcast_data_1024;
  reg [1-1:0] _eq_data_1040;
  reg [1-1:0] _eq_data_1044;
  reg [1-1:0] _eq_data_1047;
  reg [1-1:0] _eq_data_1050;
  reg [1-1:0] _eq_data_1054;
  reg [1-1:0] _eq_data_1057;
  reg [1-1:0] _eq_data_1060;
  reg [1-1:0] _eq_data_1064;
  reg [1-1:0] _eq_data_1067;
  reg [1-1:0] _eq_data_1070;
  reg [1-1:0] _eq_data_1074;
  reg [1-1:0] _eq_data_1077;
  reg [1-1:0] _eq_data_1080;
  reg [1-1:0] _eq_data_1084;
  reg [1-1:0] _eq_data_1087;
  reg [1-1:0] _eq_data_1090;
  reg [1-1:0] _eq_data_1094;
  reg [1-1:0] _eq_data_1097;
  reg [1-1:0] _eq_data_1100;
  reg [1-1:0] _eq_data_1104;
  reg [1-1:0] _eq_data_1107;
  reg [1-1:0] _eq_data_1110;
  reg [1-1:0] _eq_data_1114;
  reg [1-1:0] _eq_data_1117;
  reg [1-1:0] _eq_data_1120;
  reg [1-1:0] _eq_data_1124;
  reg [1-1:0] _eq_data_1127;
  reg [1-1:0] _eq_data_1130;
  reg [1-1:0] _eq_data_1134;
  reg [1-1:0] _eq_data_1137;
  reg [1-1:0] _eq_data_1140;
  reg [1-1:0] _eq_data_1144;
  reg [1-1:0] _eq_data_1147;
  reg [1-1:0] _eq_data_1150;
  reg [1-1:0] _eq_data_1154;
  reg [1-1:0] _eq_data_1157;
  reg [1-1:0] _eq_data_1160;
  reg [1-1:0] _eq_data_1164;
  reg [1-1:0] _eq_data_1167;
  reg [1-1:0] _eq_data_1170;
  reg [1-1:0] _eq_data_1174;
  reg [1-1:0] _eq_data_1177;
  reg [1-1:0] _eq_data_1180;
  reg [1-1:0] _eq_data_1184;
  reg [1-1:0] _eq_data_1187;
  reg [1-1:0] _eq_data_1190;
  reg [1-1:0] _eq_data_1194;
  reg [1-1:0] _eq_data_1197;
  reg [1-1:0] _eq_data_1200;
  reg [1-1:0] _eq_data_1204;
  reg [1-1:0] _eq_data_1207;
  reg [1-1:0] _eq_data_1210;
  reg [1-1:0] _eq_data_1214;
  reg [1-1:0] _eq_data_1217;
  wire [16-1:0] _slice_data_1348;
  assign _slice_data_1348 = stream_conv2d_4_source_29_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1349;
  assign _reinterpretcast_src_1349 = _slice_data_1348;
  wire signed [16-1:0] _reinterpretcast_data_1349;
  assign _reinterpretcast_data_1349 = _reinterpretcast_src_1349;
  wire [16-1:0] _slice_data_1352;
  assign _slice_data_1352 = stream_conv2d_4_source_29_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1353;
  assign _reinterpretcast_src_1353 = _slice_data_1352;
  wire signed [16-1:0] _reinterpretcast_data_1353;
  assign _reinterpretcast_data_1353 = _reinterpretcast_src_1353;
  wire [16-1:0] _slice_data_1356;
  assign _slice_data_1356 = stream_conv2d_4_source_30_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1357;
  assign _reinterpretcast_src_1357 = _slice_data_1356;
  wire signed [16-1:0] _reinterpretcast_data_1357;
  assign _reinterpretcast_data_1357 = _reinterpretcast_src_1357;
  wire [16-1:0] _slice_data_1360;
  assign _slice_data_1360 = stream_conv2d_4_source_30_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1361;
  assign _reinterpretcast_src_1361 = _slice_data_1360;
  wire signed [16-1:0] _reinterpretcast_data_1361;
  assign _reinterpretcast_data_1361 = _reinterpretcast_src_1361;
  wire [16-1:0] _slice_data_1364;
  assign _slice_data_1364 = stream_conv2d_4_source_31_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1365;
  assign _reinterpretcast_src_1365 = _slice_data_1364;
  wire signed [16-1:0] _reinterpretcast_data_1365;
  assign _reinterpretcast_data_1365 = _reinterpretcast_src_1365;
  wire [16-1:0] _slice_data_1368;
  assign _slice_data_1368 = stream_conv2d_4_source_31_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1369;
  assign _reinterpretcast_src_1369 = _slice_data_1368;
  wire signed [16-1:0] _reinterpretcast_data_1369;
  assign _reinterpretcast_data_1369 = _reinterpretcast_src_1369;
  wire [16-1:0] _slice_data_1372;
  assign _slice_data_1372 = stream_conv2d_4_source_32_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1373;
  assign _reinterpretcast_src_1373 = _slice_data_1372;
  wire signed [16-1:0] _reinterpretcast_data_1373;
  assign _reinterpretcast_data_1373 = _reinterpretcast_src_1373;
  wire [16-1:0] _slice_data_1376;
  assign _slice_data_1376 = stream_conv2d_4_source_32_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1377;
  assign _reinterpretcast_src_1377 = _slice_data_1376;
  wire signed [16-1:0] _reinterpretcast_data_1377;
  assign _reinterpretcast_data_1377 = _reinterpretcast_src_1377;
  wire [16-1:0] _slice_data_1380;
  assign _slice_data_1380 = stream_conv2d_4_source_33_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1381;
  assign _reinterpretcast_src_1381 = _slice_data_1380;
  wire signed [16-1:0] _reinterpretcast_data_1381;
  assign _reinterpretcast_data_1381 = _reinterpretcast_src_1381;
  wire [16-1:0] _slice_data_1384;
  assign _slice_data_1384 = stream_conv2d_4_source_33_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1385;
  assign _reinterpretcast_src_1385 = _slice_data_1384;
  wire signed [16-1:0] _reinterpretcast_data_1385;
  assign _reinterpretcast_data_1385 = _reinterpretcast_src_1385;
  wire [16-1:0] _slice_data_1388;
  assign _slice_data_1388 = stream_conv2d_4_source_34_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1389;
  assign _reinterpretcast_src_1389 = _slice_data_1388;
  wire signed [16-1:0] _reinterpretcast_data_1389;
  assign _reinterpretcast_data_1389 = _reinterpretcast_src_1389;
  wire [16-1:0] _slice_data_1392;
  assign _slice_data_1392 = stream_conv2d_4_source_34_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1393;
  assign _reinterpretcast_src_1393 = _slice_data_1392;
  wire signed [16-1:0] _reinterpretcast_data_1393;
  assign _reinterpretcast_data_1393 = _reinterpretcast_src_1393;
  wire [16-1:0] _slice_data_1396;
  assign _slice_data_1396 = stream_conv2d_4_source_35_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1397;
  assign _reinterpretcast_src_1397 = _slice_data_1396;
  wire signed [16-1:0] _reinterpretcast_data_1397;
  assign _reinterpretcast_data_1397 = _reinterpretcast_src_1397;
  wire [16-1:0] _slice_data_1400;
  assign _slice_data_1400 = stream_conv2d_4_source_35_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1401;
  assign _reinterpretcast_src_1401 = _slice_data_1400;
  wire signed [16-1:0] _reinterpretcast_data_1401;
  assign _reinterpretcast_data_1401 = _reinterpretcast_src_1401;
  wire [16-1:0] _slice_data_1404;
  assign _slice_data_1404 = stream_conv2d_4_source_36_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1405;
  assign _reinterpretcast_src_1405 = _slice_data_1404;
  wire signed [16-1:0] _reinterpretcast_data_1405;
  assign _reinterpretcast_data_1405 = _reinterpretcast_src_1405;
  wire [16-1:0] _slice_data_1408;
  assign _slice_data_1408 = stream_conv2d_4_source_36_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1409;
  assign _reinterpretcast_src_1409 = _slice_data_1408;
  wire signed [16-1:0] _reinterpretcast_data_1409;
  assign _reinterpretcast_data_1409 = _reinterpretcast_src_1409;
  wire [16-1:0] _slice_data_1412;
  assign _slice_data_1412 = stream_conv2d_4_source_37_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1413;
  assign _reinterpretcast_src_1413 = _slice_data_1412;
  wire signed [16-1:0] _reinterpretcast_data_1413;
  assign _reinterpretcast_data_1413 = _reinterpretcast_src_1413;
  wire [16-1:0] _slice_data_1416;
  assign _slice_data_1416 = stream_conv2d_4_source_37_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1417;
  assign _reinterpretcast_src_1417 = _slice_data_1416;
  wire signed [16-1:0] _reinterpretcast_data_1417;
  assign _reinterpretcast_data_1417 = _reinterpretcast_src_1417;
  wire [16-1:0] _slice_data_1456;
  assign _slice_data_1456 = stream_conv2d_4_source_38_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1457;
  assign _reinterpretcast_src_1457 = _slice_data_1456;
  wire signed [16-1:0] _reinterpretcast_data_1457;
  assign _reinterpretcast_data_1457 = _reinterpretcast_src_1457;
  wire [16-1:0] _slice_data_1460;
  assign _slice_data_1460 = stream_conv2d_4_source_38_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1461;
  assign _reinterpretcast_src_1461 = _slice_data_1460;
  wire signed [16-1:0] _reinterpretcast_data_1461;
  assign _reinterpretcast_data_1461 = _reinterpretcast_src_1461;
  wire [16-1:0] _slice_data_1464;
  assign _slice_data_1464 = stream_conv2d_4_source_39_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1465;
  assign _reinterpretcast_src_1465 = _slice_data_1464;
  wire signed [16-1:0] _reinterpretcast_data_1465;
  assign _reinterpretcast_data_1465 = _reinterpretcast_src_1465;
  wire [16-1:0] _slice_data_1468;
  assign _slice_data_1468 = stream_conv2d_4_source_39_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1469;
  assign _reinterpretcast_src_1469 = _slice_data_1468;
  wire signed [16-1:0] _reinterpretcast_data_1469;
  assign _reinterpretcast_data_1469 = _reinterpretcast_src_1469;
  wire [16-1:0] _slice_data_1472;
  assign _slice_data_1472 = stream_conv2d_4_source_40_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1473;
  assign _reinterpretcast_src_1473 = _slice_data_1472;
  wire signed [16-1:0] _reinterpretcast_data_1473;
  assign _reinterpretcast_data_1473 = _reinterpretcast_src_1473;
  wire [16-1:0] _slice_data_1476;
  assign _slice_data_1476 = stream_conv2d_4_source_40_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1477;
  assign _reinterpretcast_src_1477 = _slice_data_1476;
  wire signed [16-1:0] _reinterpretcast_data_1477;
  assign _reinterpretcast_data_1477 = _reinterpretcast_src_1477;
  wire [16-1:0] _slice_data_1480;
  assign _slice_data_1480 = stream_conv2d_4_source_41_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1481;
  assign _reinterpretcast_src_1481 = _slice_data_1480;
  wire signed [16-1:0] _reinterpretcast_data_1481;
  assign _reinterpretcast_data_1481 = _reinterpretcast_src_1481;
  wire [16-1:0] _slice_data_1484;
  assign _slice_data_1484 = stream_conv2d_4_source_41_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1485;
  assign _reinterpretcast_src_1485 = _slice_data_1484;
  wire signed [16-1:0] _reinterpretcast_data_1485;
  assign _reinterpretcast_data_1485 = _reinterpretcast_src_1485;
  wire [16-1:0] _slice_data_1488;
  assign _slice_data_1488 = stream_conv2d_4_source_42_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1489;
  assign _reinterpretcast_src_1489 = _slice_data_1488;
  wire signed [16-1:0] _reinterpretcast_data_1489;
  assign _reinterpretcast_data_1489 = _reinterpretcast_src_1489;
  wire [16-1:0] _slice_data_1492;
  assign _slice_data_1492 = stream_conv2d_4_source_42_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1493;
  assign _reinterpretcast_src_1493 = _slice_data_1492;
  wire signed [16-1:0] _reinterpretcast_data_1493;
  assign _reinterpretcast_data_1493 = _reinterpretcast_src_1493;
  wire [16-1:0] _slice_data_1496;
  assign _slice_data_1496 = stream_conv2d_4_source_43_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1497;
  assign _reinterpretcast_src_1497 = _slice_data_1496;
  wire signed [16-1:0] _reinterpretcast_data_1497;
  assign _reinterpretcast_data_1497 = _reinterpretcast_src_1497;
  wire [16-1:0] _slice_data_1500;
  assign _slice_data_1500 = stream_conv2d_4_source_43_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1501;
  assign _reinterpretcast_src_1501 = _slice_data_1500;
  wire signed [16-1:0] _reinterpretcast_data_1501;
  assign _reinterpretcast_data_1501 = _reinterpretcast_src_1501;
  wire [16-1:0] _slice_data_1504;
  assign _slice_data_1504 = stream_conv2d_4_source_44_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1505;
  assign _reinterpretcast_src_1505 = _slice_data_1504;
  wire signed [16-1:0] _reinterpretcast_data_1505;
  assign _reinterpretcast_data_1505 = _reinterpretcast_src_1505;
  wire [16-1:0] _slice_data_1508;
  assign _slice_data_1508 = stream_conv2d_4_source_44_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1509;
  assign _reinterpretcast_src_1509 = _slice_data_1508;
  wire signed [16-1:0] _reinterpretcast_data_1509;
  assign _reinterpretcast_data_1509 = _reinterpretcast_src_1509;
  wire [16-1:0] _slice_data_1512;
  assign _slice_data_1512 = stream_conv2d_4_source_45_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1513;
  assign _reinterpretcast_src_1513 = _slice_data_1512;
  wire signed [16-1:0] _reinterpretcast_data_1513;
  assign _reinterpretcast_data_1513 = _reinterpretcast_src_1513;
  wire [16-1:0] _slice_data_1516;
  assign _slice_data_1516 = stream_conv2d_4_source_45_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1517;
  assign _reinterpretcast_src_1517 = _slice_data_1516;
  wire signed [16-1:0] _reinterpretcast_data_1517;
  assign _reinterpretcast_data_1517 = _reinterpretcast_src_1517;
  wire [16-1:0] _slice_data_1520;
  assign _slice_data_1520 = stream_conv2d_4_source_46_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1521;
  assign _reinterpretcast_src_1521 = _slice_data_1520;
  wire signed [16-1:0] _reinterpretcast_data_1521;
  assign _reinterpretcast_data_1521 = _reinterpretcast_src_1521;
  wire [16-1:0] _slice_data_1524;
  assign _slice_data_1524 = stream_conv2d_4_source_46_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1525;
  assign _reinterpretcast_src_1525 = _slice_data_1524;
  wire signed [16-1:0] _reinterpretcast_data_1525;
  assign _reinterpretcast_data_1525 = _reinterpretcast_src_1525;
  wire [1-1:0] _pointer_data_1562;
  assign _pointer_data_1562 = stream_conv2d_4_parameter_3_data[1'sd0];
  wire [1-1:0] _pointer_data_1564;
  assign _pointer_data_1564 = stream_conv2d_4_parameter_3_data[2'sd1];
  wire [1-1:0] _pointer_data_1566;
  assign _pointer_data_1566 = stream_conv2d_4_parameter_3_data[3'sd2];
  wire [1-1:0] _pointer_data_1568;
  assign _pointer_data_1568 = stream_conv2d_4_parameter_3_data[3'sd3];
  wire [1-1:0] _pointer_data_1570;
  assign _pointer_data_1570 = stream_conv2d_4_parameter_3_data[4'sd4];
  wire [1-1:0] _pointer_data_1572;
  assign _pointer_data_1572 = stream_conv2d_4_parameter_3_data[4'sd5];
  wire [1-1:0] _pointer_data_1574;
  assign _pointer_data_1574 = stream_conv2d_4_parameter_3_data[4'sd6];
  wire [1-1:0] _pointer_data_1576;
  assign _pointer_data_1576 = stream_conv2d_4_parameter_3_data[4'sd7];
  wire [1-1:0] _pointer_data_1578;
  assign _pointer_data_1578 = stream_conv2d_4_parameter_3_data[5'sd8];
  reg [16-1:0] _plus_data_1615;
  reg [16-1:0] _plus_data_1634;
  reg [16-1:0] _plus_data_1653;
  reg [16-1:0] _plus_data_1672;
  reg [16-1:0] _plus_data_1691;
  reg [16-1:0] _plus_data_1710;
  reg [16-1:0] _plus_data_1729;
  reg [16-1:0] _plus_data_1748;
  reg [16-1:0] _plus_data_1767;
  reg [16-1:0] _plus_data_1804;
  reg [16-1:0] _plus_data_1823;
  reg [16-1:0] _plus_data_1842;
  reg [16-1:0] _plus_data_1861;
  reg [16-1:0] _plus_data_1880;
  reg [16-1:0] _plus_data_1899;
  reg [16-1:0] _plus_data_1918;
  reg [16-1:0] _plus_data_1937;
  reg [16-1:0] _plus_data_1956;
  reg [16-1:0] _plus_data_1972;
  reg [16-1:0] _plus_data_1991;
  reg [16-1:0] _plus_data_2033;
  reg [16-1:0] _plus_data_2052;
  reg [16-1:0] _plus_data_2071;
  reg [16-1:0] _plus_data_2090;
  reg [16-1:0] _plus_data_2109;
  reg [16-1:0] _plus_data_2128;
  reg [16-1:0] _plus_data_2147;
  reg [16-1:0] _plus_data_2166;
  reg [16-1:0] _plus_data_2185;
  reg [16-1:0] _plus_data_2222;
  reg [16-1:0] _plus_data_2241;
  reg [16-1:0] _plus_data_2260;
  reg [16-1:0] _plus_data_2279;
  reg [16-1:0] _plus_data_2298;
  reg [16-1:0] _plus_data_2317;
  reg [16-1:0] _plus_data_2336;
  reg [16-1:0] _plus_data_2355;
  reg [16-1:0] _plus_data_2374;
  reg [16-1:0] _plus_data_2390;
  reg [16-1:0] _plus_data_2409;
  reg [1-1:0] __delay_data_2642_pointer_955;
  reg [32-1:0] __delay_data_2644__variable_1033;
  reg [32-1:0] __delay_data_2645__variable_1032;
  reg [32-1:0] __delay_data_2646__variable_1031;
  reg [32-1:0] __delay_data_2647__variable_1036;
  reg [32-1:0] __delay_data_2648__variable_1035;
  reg [32-1:0] __delay_data_2649__variable_1034;
  reg [32-1:0] __delay_data_2650__variable_1039;
  reg [32-1:0] __delay_data_2651__variable_1038;
  reg [32-1:0] __delay_data_2652__variable_1037;
  reg [1-1:0] __delay_data_2655_pointer_1562;
  reg signed [16-1:0] __delay_data_2658_reinterpretcast_1349;
  reg [1-1:0] __delay_data_2663_pointer_961;
  reg signed [16-1:0] __delay_data_2667_reinterpretcast_1353;
  reg [1-1:0] __delay_data_2674_pointer_1564;
  reg signed [16-1:0] __delay_data_2677_reinterpretcast_1357;
  reg signed [16-1:0] __delay_data_2684_reinterpretcast_1361;
  reg [1-1:0] __delay_data_2691_pointer_1566;
  reg signed [16-1:0] __delay_data_2694_reinterpretcast_1365;
  reg signed [16-1:0] __delay_data_2701_reinterpretcast_1369;
  reg [1-1:0] __delay_data_2708_pointer_1568;
  reg signed [16-1:0] __delay_data_2711_reinterpretcast_1373;
  reg signed [16-1:0] __delay_data_2718_reinterpretcast_1377;
  reg [1-1:0] __delay_data_2725_pointer_1570;
  reg signed [16-1:0] __delay_data_2728_reinterpretcast_1381;
  reg signed [16-1:0] __delay_data_2735_reinterpretcast_1385;
  reg [1-1:0] __delay_data_2742_pointer_1572;
  reg signed [16-1:0] __delay_data_2745_reinterpretcast_1389;
  reg signed [16-1:0] __delay_data_2752_reinterpretcast_1393;
  reg [1-1:0] __delay_data_2759_pointer_1574;
  reg signed [16-1:0] __delay_data_2762_reinterpretcast_1397;
  reg signed [16-1:0] __delay_data_2769_reinterpretcast_1401;
  reg [1-1:0] __delay_data_2776_pointer_1576;
  reg signed [16-1:0] __delay_data_2779_reinterpretcast_1405;
  reg signed [16-1:0] __delay_data_2786_reinterpretcast_1409;
  reg [1-1:0] __delay_data_2793_pointer_1578;
  reg signed [16-1:0] __delay_data_2796_reinterpretcast_1413;
  reg signed [16-1:0] __delay_data_2803_reinterpretcast_1417;
  reg [1-1:0] __delay_data_2808__variable_951;
  reg [6-1:0] __delay_data_2839__variable_946;
  reg signed [16-1:0] __delay_data_2855_reinterpretcast_1457;
  reg signed [16-1:0] __delay_data_2860_reinterpretcast_1461;
  reg signed [16-1:0] __delay_data_2865_reinterpretcast_1465;
  reg signed [16-1:0] __delay_data_2870_reinterpretcast_1469;
  reg signed [16-1:0] __delay_data_2875_reinterpretcast_1473;
  reg signed [16-1:0] __delay_data_2880_reinterpretcast_1477;
  reg signed [16-1:0] __delay_data_2885_reinterpretcast_1481;
  reg signed [16-1:0] __delay_data_2890_reinterpretcast_1485;
  reg signed [16-1:0] __delay_data_2895_reinterpretcast_1489;
  reg signed [16-1:0] __delay_data_2900_reinterpretcast_1493;
  reg signed [16-1:0] __delay_data_2905_reinterpretcast_1497;
  reg signed [16-1:0] __delay_data_2910_reinterpretcast_1501;
  reg signed [16-1:0] __delay_data_2915_reinterpretcast_1505;
  reg signed [16-1:0] __delay_data_2920_reinterpretcast_1509;
  reg signed [16-1:0] __delay_data_2925_reinterpretcast_1513;
  reg signed [16-1:0] __delay_data_2930_reinterpretcast_1517;
  reg signed [16-1:0] __delay_data_2935_reinterpretcast_1521;
  reg signed [16-1:0] __delay_data_2940_reinterpretcast_1525;
  reg signed [16-1:0] __delay_data_2960_cond_978;
  reg signed [16-1:0] __delay_data_2982_cond_990;
  reg signed [16-1:0] __delay_data_3028_cond_977;
  reg signed [16-1:0] __delay_data_3050_cond_989;
  reg [1-1:0] _eq_data_959;
  reg [1-1:0] _eq_data_965;
  wire signed [32-1:0] _cond_data_1042;
  assign _cond_data_1042 = (_eq_data_1040)? __delay_data_2644__variable_1033 : 1'sd0;
  wire signed [32-1:0] _cond_data_1046;
  assign _cond_data_1046 = (_eq_data_1044)? __delay_data_2645__variable_1032 : _cond_data_1042;
  wire signed [32-1:0] _cond_data_1049;
  assign _cond_data_1049 = (_eq_data_1047)? __delay_data_2646__variable_1031 : _cond_data_1046;
  wire signed [32-1:0] _cond_data_1052;
  assign _cond_data_1052 = (_eq_data_1050)? __delay_data_2646__variable_1031 : 1'sd0;
  wire signed [32-1:0] _cond_data_1056;
  assign _cond_data_1056 = (_eq_data_1054)? __delay_data_2644__variable_1033 : _cond_data_1052;
  wire signed [32-1:0] _cond_data_1059;
  assign _cond_data_1059 = (_eq_data_1057)? __delay_data_2645__variable_1032 : _cond_data_1056;
  wire signed [32-1:0] _cond_data_1062;
  assign _cond_data_1062 = (_eq_data_1060)? __delay_data_2645__variable_1032 : 1'sd0;
  wire signed [32-1:0] _cond_data_1066;
  assign _cond_data_1066 = (_eq_data_1064)? __delay_data_2646__variable_1031 : _cond_data_1062;
  wire signed [32-1:0] _cond_data_1069;
  assign _cond_data_1069 = (_eq_data_1067)? __delay_data_2644__variable_1033 : _cond_data_1066;
  wire signed [32-1:0] _cond_data_1072;
  assign _cond_data_1072 = (_eq_data_1070)? __delay_data_2647__variable_1036 : 1'sd0;
  wire signed [32-1:0] _cond_data_1076;
  assign _cond_data_1076 = (_eq_data_1074)? __delay_data_2648__variable_1035 : _cond_data_1072;
  wire signed [32-1:0] _cond_data_1079;
  assign _cond_data_1079 = (_eq_data_1077)? __delay_data_2649__variable_1034 : _cond_data_1076;
  wire signed [32-1:0] _cond_data_1082;
  assign _cond_data_1082 = (_eq_data_1080)? __delay_data_2649__variable_1034 : 1'sd0;
  wire signed [32-1:0] _cond_data_1086;
  assign _cond_data_1086 = (_eq_data_1084)? __delay_data_2647__variable_1036 : _cond_data_1082;
  wire signed [32-1:0] _cond_data_1089;
  assign _cond_data_1089 = (_eq_data_1087)? __delay_data_2648__variable_1035 : _cond_data_1086;
  wire signed [32-1:0] _cond_data_1092;
  assign _cond_data_1092 = (_eq_data_1090)? __delay_data_2648__variable_1035 : 1'sd0;
  wire signed [32-1:0] _cond_data_1096;
  assign _cond_data_1096 = (_eq_data_1094)? __delay_data_2649__variable_1034 : _cond_data_1092;
  wire signed [32-1:0] _cond_data_1099;
  assign _cond_data_1099 = (_eq_data_1097)? __delay_data_2647__variable_1036 : _cond_data_1096;
  wire signed [32-1:0] _cond_data_1102;
  assign _cond_data_1102 = (_eq_data_1100)? __delay_data_2650__variable_1039 : 1'sd0;
  wire signed [32-1:0] _cond_data_1106;
  assign _cond_data_1106 = (_eq_data_1104)? __delay_data_2651__variable_1038 : _cond_data_1102;
  wire signed [32-1:0] _cond_data_1109;
  assign _cond_data_1109 = (_eq_data_1107)? __delay_data_2652__variable_1037 : _cond_data_1106;
  wire signed [32-1:0] _cond_data_1112;
  assign _cond_data_1112 = (_eq_data_1110)? __delay_data_2652__variable_1037 : 1'sd0;
  wire signed [32-1:0] _cond_data_1116;
  assign _cond_data_1116 = (_eq_data_1114)? __delay_data_2650__variable_1039 : _cond_data_1112;
  wire signed [32-1:0] _cond_data_1119;
  assign _cond_data_1119 = (_eq_data_1117)? __delay_data_2651__variable_1038 : _cond_data_1116;
  wire signed [32-1:0] _cond_data_1122;
  assign _cond_data_1122 = (_eq_data_1120)? __delay_data_2651__variable_1038 : 1'sd0;
  wire signed [32-1:0] _cond_data_1126;
  assign _cond_data_1126 = (_eq_data_1124)? __delay_data_2652__variable_1037 : _cond_data_1122;
  wire signed [32-1:0] _cond_data_1129;
  assign _cond_data_1129 = (_eq_data_1127)? __delay_data_2650__variable_1039 : _cond_data_1126;
  wire signed [32-1:0] _cond_data_1132;
  assign _cond_data_1132 = (_eq_data_1130)? _cond_data_1109 : 1'sd0;
  wire signed [32-1:0] _cond_data_1136;
  assign _cond_data_1136 = (_eq_data_1134)? _cond_data_1079 : _cond_data_1132;
  wire signed [32-1:0] _cond_data_1139;
  assign _cond_data_1139 = (_eq_data_1137)? _cond_data_1049 : _cond_data_1136;
  wire signed [32-1:0] _cond_data_1142;
  assign _cond_data_1142 = (_eq_data_1140)? _cond_data_1049 : 1'sd0;
  wire signed [32-1:0] _cond_data_1146;
  assign _cond_data_1146 = (_eq_data_1144)? _cond_data_1109 : _cond_data_1142;
  wire signed [32-1:0] _cond_data_1149;
  assign _cond_data_1149 = (_eq_data_1147)? _cond_data_1079 : _cond_data_1146;
  wire signed [32-1:0] _cond_data_1152;
  assign _cond_data_1152 = (_eq_data_1150)? _cond_data_1079 : 1'sd0;
  wire signed [32-1:0] _cond_data_1156;
  assign _cond_data_1156 = (_eq_data_1154)? _cond_data_1049 : _cond_data_1152;
  wire signed [32-1:0] _cond_data_1159;
  assign _cond_data_1159 = (_eq_data_1157)? _cond_data_1109 : _cond_data_1156;
  wire signed [32-1:0] _cond_data_1162;
  assign _cond_data_1162 = (_eq_data_1160)? _cond_data_1119 : 1'sd0;
  wire signed [32-1:0] _cond_data_1166;
  assign _cond_data_1166 = (_eq_data_1164)? _cond_data_1089 : _cond_data_1162;
  wire signed [32-1:0] _cond_data_1169;
  assign _cond_data_1169 = (_eq_data_1167)? _cond_data_1059 : _cond_data_1166;
  wire signed [32-1:0] _cond_data_1172;
  assign _cond_data_1172 = (_eq_data_1170)? _cond_data_1059 : 1'sd0;
  wire signed [32-1:0] _cond_data_1176;
  assign _cond_data_1176 = (_eq_data_1174)? _cond_data_1119 : _cond_data_1172;
  wire signed [32-1:0] _cond_data_1179;
  assign _cond_data_1179 = (_eq_data_1177)? _cond_data_1089 : _cond_data_1176;
  wire signed [32-1:0] _cond_data_1182;
  assign _cond_data_1182 = (_eq_data_1180)? _cond_data_1089 : 1'sd0;
  wire signed [32-1:0] _cond_data_1186;
  assign _cond_data_1186 = (_eq_data_1184)? _cond_data_1059 : _cond_data_1182;
  wire signed [32-1:0] _cond_data_1189;
  assign _cond_data_1189 = (_eq_data_1187)? _cond_data_1119 : _cond_data_1186;
  wire signed [32-1:0] _cond_data_1192;
  assign _cond_data_1192 = (_eq_data_1190)? _cond_data_1129 : 1'sd0;
  wire signed [32-1:0] _cond_data_1196;
  assign _cond_data_1196 = (_eq_data_1194)? _cond_data_1099 : _cond_data_1192;
  wire signed [32-1:0] _cond_data_1199;
  assign _cond_data_1199 = (_eq_data_1197)? _cond_data_1069 : _cond_data_1196;
  wire signed [32-1:0] _cond_data_1202;
  assign _cond_data_1202 = (_eq_data_1200)? _cond_data_1069 : 1'sd0;
  wire signed [32-1:0] _cond_data_1206;
  assign _cond_data_1206 = (_eq_data_1204)? _cond_data_1129 : _cond_data_1202;
  wire signed [32-1:0] _cond_data_1209;
  assign _cond_data_1209 = (_eq_data_1207)? _cond_data_1099 : _cond_data_1206;
  wire signed [32-1:0] _cond_data_1212;
  assign _cond_data_1212 = (_eq_data_1210)? _cond_data_1099 : 1'sd0;
  wire signed [32-1:0] _cond_data_1216;
  assign _cond_data_1216 = (_eq_data_1214)? _cond_data_1069 : _cond_data_1212;
  wire signed [32-1:0] _cond_data_1219;
  assign _cond_data_1219 = (_eq_data_1217)? _cond_data_1129 : _cond_data_1216;
  wire [16-1:0] _slice_data_1222;
  assign _slice_data_1222 = _cond_data_1139[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1223;
  assign _reinterpretcast_src_1223 = _slice_data_1222;
  wire signed [16-1:0] _reinterpretcast_data_1223;
  assign _reinterpretcast_data_1223 = _reinterpretcast_src_1223;
  wire [16-1:0] _slice_data_1226;
  assign _slice_data_1226 = _cond_data_1139[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1227;
  assign _reinterpretcast_src_1227 = _slice_data_1226;
  wire signed [16-1:0] _reinterpretcast_data_1227;
  assign _reinterpretcast_data_1227 = _reinterpretcast_src_1227;
  wire [16-1:0] _slice_data_1230;
  assign _slice_data_1230 = _cond_data_1169[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1231;
  assign _reinterpretcast_src_1231 = _slice_data_1230;
  wire signed [16-1:0] _reinterpretcast_data_1231;
  assign _reinterpretcast_data_1231 = _reinterpretcast_src_1231;
  wire [16-1:0] _slice_data_1234;
  assign _slice_data_1234 = _cond_data_1169[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1235;
  assign _reinterpretcast_src_1235 = _slice_data_1234;
  wire signed [16-1:0] _reinterpretcast_data_1235;
  assign _reinterpretcast_data_1235 = _reinterpretcast_src_1235;
  wire [16-1:0] _slice_data_1238;
  assign _slice_data_1238 = _cond_data_1199[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1239;
  assign _reinterpretcast_src_1239 = _slice_data_1238;
  wire signed [16-1:0] _reinterpretcast_data_1239;
  assign _reinterpretcast_data_1239 = _reinterpretcast_src_1239;
  wire [16-1:0] _slice_data_1242;
  assign _slice_data_1242 = _cond_data_1199[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1243;
  assign _reinterpretcast_src_1243 = _slice_data_1242;
  wire signed [16-1:0] _reinterpretcast_data_1243;
  assign _reinterpretcast_data_1243 = _reinterpretcast_src_1243;
  wire [16-1:0] _slice_data_1246;
  assign _slice_data_1246 = _cond_data_1149[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1247;
  assign _reinterpretcast_src_1247 = _slice_data_1246;
  wire signed [16-1:0] _reinterpretcast_data_1247;
  assign _reinterpretcast_data_1247 = _reinterpretcast_src_1247;
  wire [16-1:0] _slice_data_1250;
  assign _slice_data_1250 = _cond_data_1149[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1251;
  assign _reinterpretcast_src_1251 = _slice_data_1250;
  wire signed [16-1:0] _reinterpretcast_data_1251;
  assign _reinterpretcast_data_1251 = _reinterpretcast_src_1251;
  wire [16-1:0] _slice_data_1254;
  assign _slice_data_1254 = _cond_data_1179[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1255;
  assign _reinterpretcast_src_1255 = _slice_data_1254;
  wire signed [16-1:0] _reinterpretcast_data_1255;
  assign _reinterpretcast_data_1255 = _reinterpretcast_src_1255;
  wire [16-1:0] _slice_data_1258;
  assign _slice_data_1258 = _cond_data_1179[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1259;
  assign _reinterpretcast_src_1259 = _slice_data_1258;
  wire signed [16-1:0] _reinterpretcast_data_1259;
  assign _reinterpretcast_data_1259 = _reinterpretcast_src_1259;
  wire [16-1:0] _slice_data_1262;
  assign _slice_data_1262 = _cond_data_1209[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1263;
  assign _reinterpretcast_src_1263 = _slice_data_1262;
  wire signed [16-1:0] _reinterpretcast_data_1263;
  assign _reinterpretcast_data_1263 = _reinterpretcast_src_1263;
  wire [16-1:0] _slice_data_1266;
  assign _slice_data_1266 = _cond_data_1209[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1267;
  assign _reinterpretcast_src_1267 = _slice_data_1266;
  wire signed [16-1:0] _reinterpretcast_data_1267;
  assign _reinterpretcast_data_1267 = _reinterpretcast_src_1267;
  wire [16-1:0] _slice_data_1270;
  assign _slice_data_1270 = _cond_data_1159[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1271;
  assign _reinterpretcast_src_1271 = _slice_data_1270;
  wire signed [16-1:0] _reinterpretcast_data_1271;
  assign _reinterpretcast_data_1271 = _reinterpretcast_src_1271;
  wire [16-1:0] _slice_data_1274;
  assign _slice_data_1274 = _cond_data_1159[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1275;
  assign _reinterpretcast_src_1275 = _slice_data_1274;
  wire signed [16-1:0] _reinterpretcast_data_1275;
  assign _reinterpretcast_data_1275 = _reinterpretcast_src_1275;
  wire [16-1:0] _slice_data_1278;
  assign _slice_data_1278 = _cond_data_1189[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1279;
  assign _reinterpretcast_src_1279 = _slice_data_1278;
  wire signed [16-1:0] _reinterpretcast_data_1279;
  assign _reinterpretcast_data_1279 = _reinterpretcast_src_1279;
  wire [16-1:0] _slice_data_1282;
  assign _slice_data_1282 = _cond_data_1189[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1283;
  assign _reinterpretcast_src_1283 = _slice_data_1282;
  wire signed [16-1:0] _reinterpretcast_data_1283;
  assign _reinterpretcast_data_1283 = _reinterpretcast_src_1283;
  wire [16-1:0] _slice_data_1286;
  assign _slice_data_1286 = _cond_data_1219[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1287;
  assign _reinterpretcast_src_1287 = _slice_data_1286;
  wire signed [16-1:0] _reinterpretcast_data_1287;
  assign _reinterpretcast_data_1287 = _reinterpretcast_src_1287;
  wire [16-1:0] _slice_data_1290;
  assign _slice_data_1290 = _cond_data_1219[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_1291;
  assign _reinterpretcast_src_1291 = _slice_data_1290;
  wire signed [16-1:0] _reinterpretcast_data_1291;
  assign _reinterpretcast_data_1291 = _reinterpretcast_src_1291;
  reg [1-1:0] __delay_data_2643__delay_2642_pointer_955;
  reg signed [16-1:0] __delay_data_2653_reinterpretcast_1223;
  reg [1-1:0] __delay_data_2656__delay_2655_pointer_1562;
  reg signed [16-1:0] __delay_data_2659__delay_2658_reinterpretcast_1349;
  reg [16-1:0] __delay_data_2661_plus_1615;
  reg [1-1:0] __delay_data_2664__delay_2663_pointer_961;
  reg signed [16-1:0] __delay_data_2665_reinterpretcast_1227;
  reg signed [16-1:0] __delay_data_2668__delay_2667_reinterpretcast_1353;
  reg [16-1:0] __delay_data_2670_plus_1804;
  reg signed [16-1:0] __delay_data_2672_reinterpretcast_1231;
  reg [1-1:0] __delay_data_2675__delay_2674_pointer_1564;
  reg signed [16-1:0] __delay_data_2678__delay_2677_reinterpretcast_1357;
  reg [16-1:0] __delay_data_2680_plus_1634;
  reg signed [16-1:0] __delay_data_2682_reinterpretcast_1235;
  reg signed [16-1:0] __delay_data_2685__delay_2684_reinterpretcast_1361;
  reg [16-1:0] __delay_data_2687_plus_1823;
  reg signed [16-1:0] __delay_data_2689_reinterpretcast_1239;
  reg [1-1:0] __delay_data_2692__delay_2691_pointer_1566;
  reg signed [16-1:0] __delay_data_2695__delay_2694_reinterpretcast_1365;
  reg [16-1:0] __delay_data_2697_plus_1653;
  reg signed [16-1:0] __delay_data_2699_reinterpretcast_1243;
  reg signed [16-1:0] __delay_data_2702__delay_2701_reinterpretcast_1369;
  reg [16-1:0] __delay_data_2704_plus_1842;
  reg signed [16-1:0] __delay_data_2706_reinterpretcast_1247;
  reg [1-1:0] __delay_data_2709__delay_2708_pointer_1568;
  reg signed [16-1:0] __delay_data_2712__delay_2711_reinterpretcast_1373;
  reg [16-1:0] __delay_data_2714_plus_1672;
  reg signed [16-1:0] __delay_data_2716_reinterpretcast_1251;
  reg signed [16-1:0] __delay_data_2719__delay_2718_reinterpretcast_1377;
  reg [16-1:0] __delay_data_2721_plus_1861;
  reg signed [16-1:0] __delay_data_2723_reinterpretcast_1255;
  reg [1-1:0] __delay_data_2726__delay_2725_pointer_1570;
  reg signed [16-1:0] __delay_data_2729__delay_2728_reinterpretcast_1381;
  reg [16-1:0] __delay_data_2731_plus_1691;
  reg signed [16-1:0] __delay_data_2733_reinterpretcast_1259;
  reg signed [16-1:0] __delay_data_2736__delay_2735_reinterpretcast_1385;
  reg [16-1:0] __delay_data_2738_plus_1880;
  reg signed [16-1:0] __delay_data_2740_reinterpretcast_1263;
  reg [1-1:0] __delay_data_2743__delay_2742_pointer_1572;
  reg signed [16-1:0] __delay_data_2746__delay_2745_reinterpretcast_1389;
  reg [16-1:0] __delay_data_2748_plus_1710;
  reg signed [16-1:0] __delay_data_2750_reinterpretcast_1267;
  reg signed [16-1:0] __delay_data_2753__delay_2752_reinterpretcast_1393;
  reg [16-1:0] __delay_data_2755_plus_1899;
  reg signed [16-1:0] __delay_data_2757_reinterpretcast_1271;
  reg [1-1:0] __delay_data_2760__delay_2759_pointer_1574;
  reg signed [16-1:0] __delay_data_2763__delay_2762_reinterpretcast_1397;
  reg [16-1:0] __delay_data_2765_plus_1729;
  reg signed [16-1:0] __delay_data_2767_reinterpretcast_1275;
  reg signed [16-1:0] __delay_data_2770__delay_2769_reinterpretcast_1401;
  reg [16-1:0] __delay_data_2772_plus_1918;
  reg signed [16-1:0] __delay_data_2774_reinterpretcast_1279;
  reg [1-1:0] __delay_data_2777__delay_2776_pointer_1576;
  reg signed [16-1:0] __delay_data_2780__delay_2779_reinterpretcast_1405;
  reg [16-1:0] __delay_data_2782_plus_1748;
  reg signed [16-1:0] __delay_data_2784_reinterpretcast_1283;
  reg signed [16-1:0] __delay_data_2787__delay_2786_reinterpretcast_1409;
  reg [16-1:0] __delay_data_2789_plus_1937;
  reg signed [16-1:0] __delay_data_2791_reinterpretcast_1287;
  reg [1-1:0] __delay_data_2794__delay_2793_pointer_1578;
  reg signed [16-1:0] __delay_data_2797__delay_2796_reinterpretcast_1413;
  reg [16-1:0] __delay_data_2799_plus_1767;
  reg signed [16-1:0] __delay_data_2801_reinterpretcast_1291;
  reg signed [16-1:0] __delay_data_2804__delay_2803_reinterpretcast_1417;
  reg [16-1:0] __delay_data_2806_plus_1956;
  reg [1-1:0] __delay_data_2809__delay_2808__variable_951;
  reg [16-1:0] __delay_data_2824_plus_1972;
  reg [6-1:0] __delay_data_2840__delay_2839__variable_946;
  reg signed [16-1:0] __delay_data_2856__delay_2855_reinterpretcast_1457;
  reg [16-1:0] __delay_data_2858_plus_2033;
  reg signed [16-1:0] __delay_data_2861__delay_2860_reinterpretcast_1461;
  reg [16-1:0] __delay_data_2863_plus_2222;
  reg signed [16-1:0] __delay_data_2866__delay_2865_reinterpretcast_1465;
  reg [16-1:0] __delay_data_2868_plus_2052;
  reg signed [16-1:0] __delay_data_2871__delay_2870_reinterpretcast_1469;
  reg [16-1:0] __delay_data_2873_plus_2241;
  reg signed [16-1:0] __delay_data_2876__delay_2875_reinterpretcast_1473;
  reg [16-1:0] __delay_data_2878_plus_2071;
  reg signed [16-1:0] __delay_data_2881__delay_2880_reinterpretcast_1477;
  reg [16-1:0] __delay_data_2883_plus_2260;
  reg signed [16-1:0] __delay_data_2886__delay_2885_reinterpretcast_1481;
  reg [16-1:0] __delay_data_2888_plus_2090;
  reg signed [16-1:0] __delay_data_2891__delay_2890_reinterpretcast_1485;
  reg [16-1:0] __delay_data_2893_plus_2279;
  reg signed [16-1:0] __delay_data_2896__delay_2895_reinterpretcast_1489;
  reg [16-1:0] __delay_data_2898_plus_2109;
  reg signed [16-1:0] __delay_data_2901__delay_2900_reinterpretcast_1493;
  reg [16-1:0] __delay_data_2903_plus_2298;
  reg signed [16-1:0] __delay_data_2906__delay_2905_reinterpretcast_1497;
  reg [16-1:0] __delay_data_2908_plus_2128;
  reg signed [16-1:0] __delay_data_2911__delay_2910_reinterpretcast_1501;
  reg [16-1:0] __delay_data_2913_plus_2317;
  reg signed [16-1:0] __delay_data_2916__delay_2915_reinterpretcast_1505;
  reg [16-1:0] __delay_data_2918_plus_2147;
  reg signed [16-1:0] __delay_data_2921__delay_2920_reinterpretcast_1509;
  reg [16-1:0] __delay_data_2923_plus_2336;
  reg signed [16-1:0] __delay_data_2926__delay_2925_reinterpretcast_1513;
  reg [16-1:0] __delay_data_2928_plus_2166;
  reg signed [16-1:0] __delay_data_2931__delay_2930_reinterpretcast_1517;
  reg [16-1:0] __delay_data_2933_plus_2355;
  reg signed [16-1:0] __delay_data_2936__delay_2935_reinterpretcast_1521;
  reg [16-1:0] __delay_data_2938_plus_2185;
  reg signed [16-1:0] __delay_data_2941__delay_2940_reinterpretcast_1525;
  reg [16-1:0] __delay_data_2943_plus_2374;
  reg [16-1:0] __delay_data_2945_plus_2390;
  reg signed [16-1:0] __delay_data_2961__delay_2960_cond_978;
  reg signed [16-1:0] __delay_data_2983__delay_2982_cond_990;
  reg [16-1:0] __delay_data_3005_plus_2409;
  reg signed [16-1:0] __delay_data_3029__delay_3028_cond_977;
  reg signed [16-1:0] __delay_data_3051__delay_3050_cond_989;
  reg [16-1:0] __delay_data_3073_plus_1991;
  reg [1-1:0] _land_data_960;
  reg [1-1:0] _land_data_966;
  reg signed [16-1:0] __delay_data_2654__delay_2653_reinterpretcast_1223;
  reg [1-1:0] __delay_data_2657__delay_2656__delay_2655_pointer_1562;
  reg signed [16-1:0] __delay_data_2660__delay_2659__delay_2658_reinterpretcast_1349;
  reg [16-1:0] __delay_data_2662__delay_2661_plus_1615;
  reg signed [16-1:0] __delay_data_2666__delay_2665_reinterpretcast_1227;
  reg signed [16-1:0] __delay_data_2669__delay_2668__delay_2667_reinterpretcast_1353;
  reg [16-1:0] __delay_data_2671__delay_2670_plus_1804;
  reg signed [16-1:0] __delay_data_2673__delay_2672_reinterpretcast_1231;
  reg [1-1:0] __delay_data_2676__delay_2675__delay_2674_pointer_1564;
  reg signed [16-1:0] __delay_data_2679__delay_2678__delay_2677_reinterpretcast_1357;
  reg [16-1:0] __delay_data_2681__delay_2680_plus_1634;
  reg signed [16-1:0] __delay_data_2683__delay_2682_reinterpretcast_1235;
  reg signed [16-1:0] __delay_data_2686__delay_2685__delay_2684_reinterpretcast_1361;
  reg [16-1:0] __delay_data_2688__delay_2687_plus_1823;
  reg signed [16-1:0] __delay_data_2690__delay_2689_reinterpretcast_1239;
  reg [1-1:0] __delay_data_2693__delay_2692__delay_2691_pointer_1566;
  reg signed [16-1:0] __delay_data_2696__delay_2695__delay_2694_reinterpretcast_1365;
  reg [16-1:0] __delay_data_2698__delay_2697_plus_1653;
  reg signed [16-1:0] __delay_data_2700__delay_2699_reinterpretcast_1243;
  reg signed [16-1:0] __delay_data_2703__delay_2702__delay_2701_reinterpretcast_1369;
  reg [16-1:0] __delay_data_2705__delay_2704_plus_1842;
  reg signed [16-1:0] __delay_data_2707__delay_2706_reinterpretcast_1247;
  reg [1-1:0] __delay_data_2710__delay_2709__delay_2708_pointer_1568;
  reg signed [16-1:0] __delay_data_2713__delay_2712__delay_2711_reinterpretcast_1373;
  reg [16-1:0] __delay_data_2715__delay_2714_plus_1672;
  reg signed [16-1:0] __delay_data_2717__delay_2716_reinterpretcast_1251;
  reg signed [16-1:0] __delay_data_2720__delay_2719__delay_2718_reinterpretcast_1377;
  reg [16-1:0] __delay_data_2722__delay_2721_plus_1861;
  reg signed [16-1:0] __delay_data_2724__delay_2723_reinterpretcast_1255;
  reg [1-1:0] __delay_data_2727__delay_2726__delay_2725_pointer_1570;
  reg signed [16-1:0] __delay_data_2730__delay_2729__delay_2728_reinterpretcast_1381;
  reg [16-1:0] __delay_data_2732__delay_2731_plus_1691;
  reg signed [16-1:0] __delay_data_2734__delay_2733_reinterpretcast_1259;
  reg signed [16-1:0] __delay_data_2737__delay_2736__delay_2735_reinterpretcast_1385;
  reg [16-1:0] __delay_data_2739__delay_2738_plus_1880;
  reg signed [16-1:0] __delay_data_2741__delay_2740_reinterpretcast_1263;
  reg [1-1:0] __delay_data_2744__delay_2743__delay_2742_pointer_1572;
  reg signed [16-1:0] __delay_data_2747__delay_2746__delay_2745_reinterpretcast_1389;
  reg [16-1:0] __delay_data_2749__delay_2748_plus_1710;
  reg signed [16-1:0] __delay_data_2751__delay_2750_reinterpretcast_1267;
  reg signed [16-1:0] __delay_data_2754__delay_2753__delay_2752_reinterpretcast_1393;
  reg [16-1:0] __delay_data_2756__delay_2755_plus_1899;
  reg signed [16-1:0] __delay_data_2758__delay_2757_reinterpretcast_1271;
  reg [1-1:0] __delay_data_2761__delay_2760__delay_2759_pointer_1574;
  reg signed [16-1:0] __delay_data_2764__delay_2763__delay_2762_reinterpretcast_1397;
  reg [16-1:0] __delay_data_2766__delay_2765_plus_1729;
  reg signed [16-1:0] __delay_data_2768__delay_2767_reinterpretcast_1275;
  reg signed [16-1:0] __delay_data_2771__delay_2770__delay_2769_reinterpretcast_1401;
  reg [16-1:0] __delay_data_2773__delay_2772_plus_1918;
  reg signed [16-1:0] __delay_data_2775__delay_2774_reinterpretcast_1279;
  reg [1-1:0] __delay_data_2778__delay_2777__delay_2776_pointer_1576;
  reg signed [16-1:0] __delay_data_2781__delay_2780__delay_2779_reinterpretcast_1405;
  reg [16-1:0] __delay_data_2783__delay_2782_plus_1748;
  reg signed [16-1:0] __delay_data_2785__delay_2784_reinterpretcast_1283;
  reg signed [16-1:0] __delay_data_2788__delay_2787__delay_2786_reinterpretcast_1409;
  reg [16-1:0] __delay_data_2790__delay_2789_plus_1937;
  reg signed [16-1:0] __delay_data_2792__delay_2791_reinterpretcast_1287;
  reg [1-1:0] __delay_data_2795__delay_2794__delay_2793_pointer_1578;
  reg signed [16-1:0] __delay_data_2798__delay_2797__delay_2796_reinterpretcast_1413;
  reg [16-1:0] __delay_data_2800__delay_2799_plus_1767;
  reg signed [16-1:0] __delay_data_2802__delay_2801_reinterpretcast_1291;
  reg signed [16-1:0] __delay_data_2805__delay_2804__delay_2803_reinterpretcast_1417;
  reg [16-1:0] __delay_data_2807__delay_2806_plus_1956;
  reg [1-1:0] __delay_data_2810__delay_2809__delay_2808__variable_951;
  reg [16-1:0] __delay_data_2825__delay_2824_plus_1972;
  reg [6-1:0] __delay_data_2841__delay_2840__delay_2839__variable_946;
  reg signed [16-1:0] __delay_data_2857__delay_2856__delay_2855_reinterpretcast_1457;
  reg [16-1:0] __delay_data_2859__delay_2858_plus_2033;
  reg signed [16-1:0] __delay_data_2862__delay_2861__delay_2860_reinterpretcast_1461;
  reg [16-1:0] __delay_data_2864__delay_2863_plus_2222;
  reg signed [16-1:0] __delay_data_2867__delay_2866__delay_2865_reinterpretcast_1465;
  reg [16-1:0] __delay_data_2869__delay_2868_plus_2052;
  reg signed [16-1:0] __delay_data_2872__delay_2871__delay_2870_reinterpretcast_1469;
  reg [16-1:0] __delay_data_2874__delay_2873_plus_2241;
  reg signed [16-1:0] __delay_data_2877__delay_2876__delay_2875_reinterpretcast_1473;
  reg [16-1:0] __delay_data_2879__delay_2878_plus_2071;
  reg signed [16-1:0] __delay_data_2882__delay_2881__delay_2880_reinterpretcast_1477;
  reg [16-1:0] __delay_data_2884__delay_2883_plus_2260;
  reg signed [16-1:0] __delay_data_2887__delay_2886__delay_2885_reinterpretcast_1481;
  reg [16-1:0] __delay_data_2889__delay_2888_plus_2090;
  reg signed [16-1:0] __delay_data_2892__delay_2891__delay_2890_reinterpretcast_1485;
  reg [16-1:0] __delay_data_2894__delay_2893_plus_2279;
  reg signed [16-1:0] __delay_data_2897__delay_2896__delay_2895_reinterpretcast_1489;
  reg [16-1:0] __delay_data_2899__delay_2898_plus_2109;
  reg signed [16-1:0] __delay_data_2902__delay_2901__delay_2900_reinterpretcast_1493;
  reg [16-1:0] __delay_data_2904__delay_2903_plus_2298;
  reg signed [16-1:0] __delay_data_2907__delay_2906__delay_2905_reinterpretcast_1497;
  reg [16-1:0] __delay_data_2909__delay_2908_plus_2128;
  reg signed [16-1:0] __delay_data_2912__delay_2911__delay_2910_reinterpretcast_1501;
  reg [16-1:0] __delay_data_2914__delay_2913_plus_2317;
  reg signed [16-1:0] __delay_data_2917__delay_2916__delay_2915_reinterpretcast_1505;
  reg [16-1:0] __delay_data_2919__delay_2918_plus_2147;
  reg signed [16-1:0] __delay_data_2922__delay_2921__delay_2920_reinterpretcast_1509;
  reg [16-1:0] __delay_data_2924__delay_2923_plus_2336;
  reg signed [16-1:0] __delay_data_2927__delay_2926__delay_2925_reinterpretcast_1513;
  reg [16-1:0] __delay_data_2929__delay_2928_plus_2166;
  reg signed [16-1:0] __delay_data_2932__delay_2931__delay_2930_reinterpretcast_1517;
  reg [16-1:0] __delay_data_2934__delay_2933_plus_2355;
  reg signed [16-1:0] __delay_data_2937__delay_2936__delay_2935_reinterpretcast_1521;
  reg [16-1:0] __delay_data_2939__delay_2938_plus_2185;
  reg signed [16-1:0] __delay_data_2942__delay_2941__delay_2940_reinterpretcast_1525;
  reg [16-1:0] __delay_data_2944__delay_2943_plus_2374;
  reg [16-1:0] __delay_data_2946__delay_2945_plus_2390;
  reg signed [16-1:0] __delay_data_2962__delay_2961__delay_2960_cond_978;
  reg signed [16-1:0] __delay_data_2984__delay_2983__delay_2982_cond_990;
  reg [16-1:0] __delay_data_3006__delay_3005_plus_2409;
  reg signed [16-1:0] __delay_data_3030__delay_3029__delay_3028_cond_977;
  reg signed [16-1:0] __delay_data_3052__delay_3051__delay_3050_cond_989;
  reg [16-1:0] __delay_data_3074__delay_3073_plus_1991;
  wire signed [16-1:0] _cond_data_1293;
  assign _cond_data_1293 = (_land_data_960)? 1'sd0 : __delay_data_2654__delay_2653_reinterpretcast_1223;
  wire signed [16-1:0] _cond_data_1295;
  assign _cond_data_1295 = (_land_data_960)? 1'sd0 : __delay_data_2673__delay_2672_reinterpretcast_1231;
  wire signed [16-1:0] _cond_data_1297;
  assign _cond_data_1297 = (_land_data_960)? 1'sd0 : __delay_data_2690__delay_2689_reinterpretcast_1239;
  wire signed [16-1:0] _cond_data_1299;
  assign _cond_data_1299 = (_land_data_960)? 1'sd0 : __delay_data_2707__delay_2706_reinterpretcast_1247;
  wire signed [16-1:0] _cond_data_1301;
  assign _cond_data_1301 = (_land_data_960)? 1'sd0 : __delay_data_2724__delay_2723_reinterpretcast_1255;
  wire signed [16-1:0] _cond_data_1303;
  assign _cond_data_1303 = (_land_data_960)? 1'sd0 : __delay_data_2741__delay_2740_reinterpretcast_1263;
  wire signed [16-1:0] _cond_data_1305;
  assign _cond_data_1305 = (_land_data_960)? 1'sd0 : __delay_data_2758__delay_2757_reinterpretcast_1271;
  wire signed [16-1:0] _cond_data_1307;
  assign _cond_data_1307 = (_land_data_960)? 1'sd0 : __delay_data_2775__delay_2774_reinterpretcast_1279;
  wire signed [16-1:0] _cond_data_1309;
  assign _cond_data_1309 = (_land_data_960)? 1'sd0 : __delay_data_2792__delay_2791_reinterpretcast_1287;
  wire signed [16-1:0] _cond_data_1311;
  assign _cond_data_1311 = (_land_data_966)? 1'sd0 : __delay_data_2666__delay_2665_reinterpretcast_1227;
  wire signed [16-1:0] _cond_data_1313;
  assign _cond_data_1313 = (_land_data_966)? 1'sd0 : __delay_data_2683__delay_2682_reinterpretcast_1235;
  wire signed [16-1:0] _cond_data_1315;
  assign _cond_data_1315 = (_land_data_966)? 1'sd0 : __delay_data_2700__delay_2699_reinterpretcast_1243;
  wire signed [16-1:0] _cond_data_1317;
  assign _cond_data_1317 = (_land_data_966)? 1'sd0 : __delay_data_2717__delay_2716_reinterpretcast_1251;
  wire signed [16-1:0] _cond_data_1319;
  assign _cond_data_1319 = (_land_data_966)? 1'sd0 : __delay_data_2734__delay_2733_reinterpretcast_1259;
  wire signed [16-1:0] _cond_data_1321;
  assign _cond_data_1321 = (_land_data_966)? 1'sd0 : __delay_data_2751__delay_2750_reinterpretcast_1267;
  wire signed [16-1:0] _cond_data_1323;
  assign _cond_data_1323 = (_land_data_966)? 1'sd0 : __delay_data_2768__delay_2767_reinterpretcast_1275;
  wire signed [16-1:0] _cond_data_1325;
  assign _cond_data_1325 = (_land_data_966)? 1'sd0 : __delay_data_2785__delay_2784_reinterpretcast_1283;
  wire signed [16-1:0] _cond_data_1327;
  assign _cond_data_1327 = (_land_data_966)? 1'sd0 : __delay_data_2802__delay_2801_reinterpretcast_1291;
  wire signed [16-1:0] _cond_data_1419;
  assign _cond_data_1419 = (_land_data_960)? 1'sd0 : __delay_data_2660__delay_2659__delay_2658_reinterpretcast_1349;
  wire signed [16-1:0] _cond_data_1421;
  assign _cond_data_1421 = (_land_data_960)? 1'sd0 : __delay_data_2679__delay_2678__delay_2677_reinterpretcast_1357;
  wire signed [16-1:0] _cond_data_1423;
  assign _cond_data_1423 = (_land_data_960)? 1'sd0 : __delay_data_2696__delay_2695__delay_2694_reinterpretcast_1365;
  wire signed [16-1:0] _cond_data_1425;
  assign _cond_data_1425 = (_land_data_960)? 1'sd0 : __delay_data_2713__delay_2712__delay_2711_reinterpretcast_1373;
  wire signed [16-1:0] _cond_data_1427;
  assign _cond_data_1427 = (_land_data_960)? 1'sd0 : __delay_data_2730__delay_2729__delay_2728_reinterpretcast_1381;
  wire signed [16-1:0] _cond_data_1429;
  assign _cond_data_1429 = (_land_data_960)? 1'sd0 : __delay_data_2747__delay_2746__delay_2745_reinterpretcast_1389;
  wire signed [16-1:0] _cond_data_1431;
  assign _cond_data_1431 = (_land_data_960)? 1'sd0 : __delay_data_2764__delay_2763__delay_2762_reinterpretcast_1397;
  wire signed [16-1:0] _cond_data_1433;
  assign _cond_data_1433 = (_land_data_960)? 1'sd0 : __delay_data_2781__delay_2780__delay_2779_reinterpretcast_1405;
  wire signed [16-1:0] _cond_data_1435;
  assign _cond_data_1435 = (_land_data_960)? 1'sd0 : __delay_data_2798__delay_2797__delay_2796_reinterpretcast_1413;
  wire signed [16-1:0] _cond_data_1437;
  assign _cond_data_1437 = (_land_data_966)? 1'sd0 : __delay_data_2669__delay_2668__delay_2667_reinterpretcast_1353;
  wire signed [16-1:0] _cond_data_1439;
  assign _cond_data_1439 = (_land_data_966)? 1'sd0 : __delay_data_2686__delay_2685__delay_2684_reinterpretcast_1361;
  wire signed [16-1:0] _cond_data_1441;
  assign _cond_data_1441 = (_land_data_966)? 1'sd0 : __delay_data_2703__delay_2702__delay_2701_reinterpretcast_1369;
  wire signed [16-1:0] _cond_data_1443;
  assign _cond_data_1443 = (_land_data_966)? 1'sd0 : __delay_data_2720__delay_2719__delay_2718_reinterpretcast_1377;
  wire signed [16-1:0] _cond_data_1445;
  assign _cond_data_1445 = (_land_data_966)? 1'sd0 : __delay_data_2737__delay_2736__delay_2735_reinterpretcast_1385;
  wire signed [16-1:0] _cond_data_1447;
  assign _cond_data_1447 = (_land_data_966)? 1'sd0 : __delay_data_2754__delay_2753__delay_2752_reinterpretcast_1393;
  wire signed [16-1:0] _cond_data_1449;
  assign _cond_data_1449 = (_land_data_966)? 1'sd0 : __delay_data_2771__delay_2770__delay_2769_reinterpretcast_1401;
  wire signed [16-1:0] _cond_data_1451;
  assign _cond_data_1451 = (_land_data_966)? 1'sd0 : __delay_data_2788__delay_2787__delay_2786_reinterpretcast_1409;
  wire signed [16-1:0] _cond_data_1453;
  assign _cond_data_1453 = (_land_data_966)? 1'sd0 : __delay_data_2805__delay_2804__delay_2803_reinterpretcast_1417;
  wire signed [16-1:0] _cond_data_1527;
  assign _cond_data_1527 = (_land_data_960)? 1'sd0 : __delay_data_2857__delay_2856__delay_2855_reinterpretcast_1457;
  wire signed [16-1:0] _cond_data_1529;
  assign _cond_data_1529 = (_land_data_960)? 1'sd0 : __delay_data_2867__delay_2866__delay_2865_reinterpretcast_1465;
  wire signed [16-1:0] _cond_data_1531;
  assign _cond_data_1531 = (_land_data_960)? 1'sd0 : __delay_data_2877__delay_2876__delay_2875_reinterpretcast_1473;
  wire signed [16-1:0] _cond_data_1533;
  assign _cond_data_1533 = (_land_data_960)? 1'sd0 : __delay_data_2887__delay_2886__delay_2885_reinterpretcast_1481;
  wire signed [16-1:0] _cond_data_1535;
  assign _cond_data_1535 = (_land_data_960)? 1'sd0 : __delay_data_2897__delay_2896__delay_2895_reinterpretcast_1489;
  wire signed [16-1:0] _cond_data_1537;
  assign _cond_data_1537 = (_land_data_960)? 1'sd0 : __delay_data_2907__delay_2906__delay_2905_reinterpretcast_1497;
  wire signed [16-1:0] _cond_data_1539;
  assign _cond_data_1539 = (_land_data_960)? 1'sd0 : __delay_data_2917__delay_2916__delay_2915_reinterpretcast_1505;
  wire signed [16-1:0] _cond_data_1541;
  assign _cond_data_1541 = (_land_data_960)? 1'sd0 : __delay_data_2927__delay_2926__delay_2925_reinterpretcast_1513;
  wire signed [16-1:0] _cond_data_1543;
  assign _cond_data_1543 = (_land_data_960)? 1'sd0 : __delay_data_2937__delay_2936__delay_2935_reinterpretcast_1521;
  wire signed [16-1:0] _cond_data_1545;
  assign _cond_data_1545 = (_land_data_966)? 1'sd0 : __delay_data_2862__delay_2861__delay_2860_reinterpretcast_1461;
  wire signed [16-1:0] _cond_data_1547;
  assign _cond_data_1547 = (_land_data_966)? 1'sd0 : __delay_data_2872__delay_2871__delay_2870_reinterpretcast_1469;
  wire signed [16-1:0] _cond_data_1549;
  assign _cond_data_1549 = (_land_data_966)? 1'sd0 : __delay_data_2882__delay_2881__delay_2880_reinterpretcast_1477;
  wire signed [16-1:0] _cond_data_1551;
  assign _cond_data_1551 = (_land_data_966)? 1'sd0 : __delay_data_2892__delay_2891__delay_2890_reinterpretcast_1485;
  wire signed [16-1:0] _cond_data_1553;
  assign _cond_data_1553 = (_land_data_966)? 1'sd0 : __delay_data_2902__delay_2901__delay_2900_reinterpretcast_1493;
  wire signed [16-1:0] _cond_data_1555;
  assign _cond_data_1555 = (_land_data_966)? 1'sd0 : __delay_data_2912__delay_2911__delay_2910_reinterpretcast_1501;
  wire signed [16-1:0] _cond_data_1557;
  assign _cond_data_1557 = (_land_data_966)? 1'sd0 : __delay_data_2922__delay_2921__delay_2920_reinterpretcast_1509;
  wire signed [16-1:0] _cond_data_1559;
  assign _cond_data_1559 = (_land_data_966)? 1'sd0 : __delay_data_2932__delay_2931__delay_2930_reinterpretcast_1517;
  wire signed [16-1:0] _cond_data_1561;
  assign _cond_data_1561 = (_land_data_966)? 1'sd0 : __delay_data_2942__delay_2941__delay_2940_reinterpretcast_1525;
  wire signed [16-1:0] _cond_data_1581;
  assign _cond_data_1581 = (__delay_data_2657__delay_2656__delay_2655_pointer_1562)? 1'sd0 : _cond_data_1293;
  wire signed [16-1:0] _cond_data_1583;
  assign _cond_data_1583 = (__delay_data_2676__delay_2675__delay_2674_pointer_1564)? 1'sd0 : _cond_data_1295;
  wire signed [16-1:0] _cond_data_1585;
  assign _cond_data_1585 = (__delay_data_2693__delay_2692__delay_2691_pointer_1566)? 1'sd0 : _cond_data_1297;
  wire signed [16-1:0] _cond_data_1587;
  assign _cond_data_1587 = (__delay_data_2710__delay_2709__delay_2708_pointer_1568)? 1'sd0 : _cond_data_1299;
  wire signed [16-1:0] _cond_data_1589;
  assign _cond_data_1589 = (__delay_data_2727__delay_2726__delay_2725_pointer_1570)? 1'sd0 : _cond_data_1301;
  wire signed [16-1:0] _cond_data_1591;
  assign _cond_data_1591 = (__delay_data_2744__delay_2743__delay_2742_pointer_1572)? 1'sd0 : _cond_data_1303;
  wire signed [16-1:0] _cond_data_1593;
  assign _cond_data_1593 = (__delay_data_2761__delay_2760__delay_2759_pointer_1574)? 1'sd0 : _cond_data_1305;
  wire signed [16-1:0] _cond_data_1595;
  assign _cond_data_1595 = (__delay_data_2778__delay_2777__delay_2776_pointer_1576)? 1'sd0 : _cond_data_1307;
  wire signed [16-1:0] _cond_data_1597;
  assign _cond_data_1597 = (__delay_data_2795__delay_2794__delay_2793_pointer_1578)? 1'sd0 : _cond_data_1309;
  reg signed [16-1:0] __variable_wdata_176;
  assign mul_8_x_data = __variable_wdata_176;
  reg signed [16-1:0] __variable_wdata_177;
  assign mul_8_y_data = __variable_wdata_177;
  reg [5-1:0] __variable_wdata_178;
  assign mul_8_rshift_data = __variable_wdata_178;
  reg signed [16-1:0] __variable_wdata_197;
  assign mul_9_x_data = __variable_wdata_197;
  reg signed [16-1:0] __variable_wdata_198;
  assign mul_9_y_data = __variable_wdata_198;
  reg [5-1:0] __variable_wdata_199;
  assign mul_9_rshift_data = __variable_wdata_199;
  reg signed [16-1:0] __variable_wdata_218;
  assign mul_10_x_data = __variable_wdata_218;
  reg signed [16-1:0] __variable_wdata_219;
  assign mul_10_y_data = __variable_wdata_219;
  reg [5-1:0] __variable_wdata_220;
  assign mul_10_rshift_data = __variable_wdata_220;
  reg signed [16-1:0] __variable_wdata_239;
  assign mul_11_x_data = __variable_wdata_239;
  reg signed [16-1:0] __variable_wdata_240;
  assign mul_11_y_data = __variable_wdata_240;
  reg [5-1:0] __variable_wdata_241;
  assign mul_11_rshift_data = __variable_wdata_241;
  reg signed [16-1:0] __variable_wdata_260;
  assign mul_12_x_data = __variable_wdata_260;
  reg signed [16-1:0] __variable_wdata_261;
  assign mul_12_y_data = __variable_wdata_261;
  reg [5-1:0] __variable_wdata_262;
  assign mul_12_rshift_data = __variable_wdata_262;
  assign _mul_12_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_12_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_12_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_281;
  assign mul_13_x_data = __variable_wdata_281;
  reg signed [16-1:0] __variable_wdata_282;
  assign mul_13_y_data = __variable_wdata_282;
  reg [5-1:0] __variable_wdata_283;
  assign mul_13_rshift_data = __variable_wdata_283;
  assign _mul_13_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_13_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_13_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_302;
  assign mul_14_x_data = __variable_wdata_302;
  reg signed [16-1:0] __variable_wdata_303;
  assign mul_14_y_data = __variable_wdata_303;
  reg [5-1:0] __variable_wdata_304;
  assign mul_14_rshift_data = __variable_wdata_304;
  assign _mul_14_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_14_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_14_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_323;
  assign mul_15_x_data = __variable_wdata_323;
  reg signed [16-1:0] __variable_wdata_324;
  assign mul_15_y_data = __variable_wdata_324;
  reg [5-1:0] __variable_wdata_325;
  assign mul_15_rshift_data = __variable_wdata_325;
  assign _mul_15_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_15_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_15_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_344;
  assign mul_16_x_data = __variable_wdata_344;
  reg signed [16-1:0] __variable_wdata_345;
  assign mul_16_y_data = __variable_wdata_345;
  reg [5-1:0] __variable_wdata_346;
  assign mul_16_rshift_data = __variable_wdata_346;
  assign _mul_16_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_16_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_16_stream_internal_oready;
  wire signed [16-1:0] _cond_data_1770;
  assign _cond_data_1770 = (__delay_data_2657__delay_2656__delay_2655_pointer_1562)? 1'sd0 : _cond_data_1311;
  wire signed [16-1:0] _cond_data_1772;
  assign _cond_data_1772 = (__delay_data_2676__delay_2675__delay_2674_pointer_1564)? 1'sd0 : _cond_data_1313;
  wire signed [16-1:0] _cond_data_1774;
  assign _cond_data_1774 = (__delay_data_2693__delay_2692__delay_2691_pointer_1566)? 1'sd0 : _cond_data_1315;
  wire signed [16-1:0] _cond_data_1776;
  assign _cond_data_1776 = (__delay_data_2710__delay_2709__delay_2708_pointer_1568)? 1'sd0 : _cond_data_1317;
  wire signed [16-1:0] _cond_data_1778;
  assign _cond_data_1778 = (__delay_data_2727__delay_2726__delay_2725_pointer_1570)? 1'sd0 : _cond_data_1319;
  wire signed [16-1:0] _cond_data_1780;
  assign _cond_data_1780 = (__delay_data_2744__delay_2743__delay_2742_pointer_1572)? 1'sd0 : _cond_data_1321;
  wire signed [16-1:0] _cond_data_1782;
  assign _cond_data_1782 = (__delay_data_2761__delay_2760__delay_2759_pointer_1574)? 1'sd0 : _cond_data_1323;
  wire signed [16-1:0] _cond_data_1784;
  assign _cond_data_1784 = (__delay_data_2778__delay_2777__delay_2776_pointer_1576)? 1'sd0 : _cond_data_1325;
  wire signed [16-1:0] _cond_data_1786;
  assign _cond_data_1786 = (__delay_data_2795__delay_2794__delay_2793_pointer_1578)? 1'sd0 : _cond_data_1327;
  reg signed [16-1:0] __variable_wdata_365;
  assign mul_17_x_data = __variable_wdata_365;
  reg signed [16-1:0] __variable_wdata_366;
  assign mul_17_y_data = __variable_wdata_366;
  reg [5-1:0] __variable_wdata_367;
  assign mul_17_rshift_data = __variable_wdata_367;
  assign _mul_17_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_17_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_17_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_386;
  assign mul_18_x_data = __variable_wdata_386;
  reg signed [16-1:0] __variable_wdata_387;
  assign mul_18_y_data = __variable_wdata_387;
  reg [5-1:0] __variable_wdata_388;
  assign mul_18_rshift_data = __variable_wdata_388;
  assign _mul_18_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_18_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_18_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_407;
  assign mul_19_x_data = __variable_wdata_407;
  reg signed [16-1:0] __variable_wdata_408;
  assign mul_19_y_data = __variable_wdata_408;
  reg [5-1:0] __variable_wdata_409;
  assign mul_19_rshift_data = __variable_wdata_409;
  assign _mul_19_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_19_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_19_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_428;
  assign mul_20_x_data = __variable_wdata_428;
  reg signed [16-1:0] __variable_wdata_429;
  assign mul_20_y_data = __variable_wdata_429;
  reg [5-1:0] __variable_wdata_430;
  assign mul_20_rshift_data = __variable_wdata_430;
  assign _mul_20_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_20_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_20_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_449;
  assign mul_21_x_data = __variable_wdata_449;
  reg signed [16-1:0] __variable_wdata_450;
  assign mul_21_y_data = __variable_wdata_450;
  reg [5-1:0] __variable_wdata_451;
  assign mul_21_rshift_data = __variable_wdata_451;
  assign _mul_21_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_21_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_21_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_470;
  assign mul_22_x_data = __variable_wdata_470;
  reg signed [16-1:0] __variable_wdata_471;
  assign mul_22_y_data = __variable_wdata_471;
  reg [5-1:0] __variable_wdata_472;
  assign mul_22_rshift_data = __variable_wdata_472;
  assign _mul_22_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_22_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_22_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_491;
  assign mul_23_x_data = __variable_wdata_491;
  reg signed [16-1:0] __variable_wdata_492;
  assign mul_23_y_data = __variable_wdata_492;
  reg [5-1:0] __variable_wdata_493;
  assign mul_23_rshift_data = __variable_wdata_493;
  assign _mul_23_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_23_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_23_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_512;
  assign mul_24_x_data = __variable_wdata_512;
  reg signed [16-1:0] __variable_wdata_513;
  assign mul_24_y_data = __variable_wdata_513;
  reg [5-1:0] __variable_wdata_514;
  assign mul_24_rshift_data = __variable_wdata_514;
  assign _mul_24_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_24_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_24_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_533;
  assign mul_25_x_data = __variable_wdata_533;
  reg signed [16-1:0] __variable_wdata_534;
  assign mul_25_y_data = __variable_wdata_534;
  reg [5-1:0] __variable_wdata_535;
  assign mul_25_rshift_data = __variable_wdata_535;
  assign _mul_25_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_25_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_25_stream_internal_oready;
  wire signed [16-1:0] _cond_data_1999;
  assign _cond_data_1999 = (__delay_data_2657__delay_2656__delay_2655_pointer_1562)? 1'sd0 : _cond_data_1293;
  wire signed [16-1:0] _cond_data_2001;
  assign _cond_data_2001 = (__delay_data_2676__delay_2675__delay_2674_pointer_1564)? 1'sd0 : _cond_data_1295;
  wire signed [16-1:0] _cond_data_2003;
  assign _cond_data_2003 = (__delay_data_2693__delay_2692__delay_2691_pointer_1566)? 1'sd0 : _cond_data_1297;
  wire signed [16-1:0] _cond_data_2005;
  assign _cond_data_2005 = (__delay_data_2710__delay_2709__delay_2708_pointer_1568)? 1'sd0 : _cond_data_1299;
  wire signed [16-1:0] _cond_data_2007;
  assign _cond_data_2007 = (__delay_data_2727__delay_2726__delay_2725_pointer_1570)? 1'sd0 : _cond_data_1301;
  wire signed [16-1:0] _cond_data_2009;
  assign _cond_data_2009 = (__delay_data_2744__delay_2743__delay_2742_pointer_1572)? 1'sd0 : _cond_data_1303;
  wire signed [16-1:0] _cond_data_2011;
  assign _cond_data_2011 = (__delay_data_2761__delay_2760__delay_2759_pointer_1574)? 1'sd0 : _cond_data_1305;
  wire signed [16-1:0] _cond_data_2013;
  assign _cond_data_2013 = (__delay_data_2778__delay_2777__delay_2776_pointer_1576)? 1'sd0 : _cond_data_1307;
  wire signed [16-1:0] _cond_data_2015;
  assign _cond_data_2015 = (__delay_data_2795__delay_2794__delay_2793_pointer_1578)? 1'sd0 : _cond_data_1309;
  reg signed [16-1:0] __variable_wdata_554;
  assign mul_26_x_data = __variable_wdata_554;
  reg signed [16-1:0] __variable_wdata_555;
  assign mul_26_y_data = __variable_wdata_555;
  reg [5-1:0] __variable_wdata_556;
  assign mul_26_rshift_data = __variable_wdata_556;
  assign _mul_26_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_26_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_26_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_575;
  assign mul_27_x_data = __variable_wdata_575;
  reg signed [16-1:0] __variable_wdata_576;
  assign mul_27_y_data = __variable_wdata_576;
  reg [5-1:0] __variable_wdata_577;
  assign mul_27_rshift_data = __variable_wdata_577;
  assign _mul_27_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_27_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_27_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_596;
  assign mul_28_x_data = __variable_wdata_596;
  reg signed [16-1:0] __variable_wdata_597;
  assign mul_28_y_data = __variable_wdata_597;
  reg [5-1:0] __variable_wdata_598;
  assign mul_28_rshift_data = __variable_wdata_598;
  assign _mul_28_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_28_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_28_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_617;
  assign mul_29_x_data = __variable_wdata_617;
  reg signed [16-1:0] __variable_wdata_618;
  assign mul_29_y_data = __variable_wdata_618;
  reg [5-1:0] __variable_wdata_619;
  assign mul_29_rshift_data = __variable_wdata_619;
  assign _mul_29_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_29_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_29_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_638;
  assign mul_30_x_data = __variable_wdata_638;
  reg signed [16-1:0] __variable_wdata_639;
  assign mul_30_y_data = __variable_wdata_639;
  reg [5-1:0] __variable_wdata_640;
  assign mul_30_rshift_data = __variable_wdata_640;
  assign _mul_30_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_30_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_30_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_659;
  assign mul_31_x_data = __variable_wdata_659;
  reg signed [16-1:0] __variable_wdata_660;
  assign mul_31_y_data = __variable_wdata_660;
  reg [5-1:0] __variable_wdata_661;
  assign mul_31_rshift_data = __variable_wdata_661;
  assign _mul_31_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_31_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_31_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_680;
  assign mul_32_x_data = __variable_wdata_680;
  reg signed [16-1:0] __variable_wdata_681;
  assign mul_32_y_data = __variable_wdata_681;
  reg [5-1:0] __variable_wdata_682;
  assign mul_32_rshift_data = __variable_wdata_682;
  assign _mul_32_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_32_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_32_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_701;
  assign mul_33_x_data = __variable_wdata_701;
  reg signed [16-1:0] __variable_wdata_702;
  assign mul_33_y_data = __variable_wdata_702;
  reg [5-1:0] __variable_wdata_703;
  assign mul_33_rshift_data = __variable_wdata_703;
  assign _mul_33_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_33_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_33_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_722;
  assign mul_34_x_data = __variable_wdata_722;
  reg signed [16-1:0] __variable_wdata_723;
  assign mul_34_y_data = __variable_wdata_723;
  reg [5-1:0] __variable_wdata_724;
  assign mul_34_rshift_data = __variable_wdata_724;
  assign _mul_34_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_34_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_34_stream_internal_oready;
  wire signed [16-1:0] _cond_data_2188;
  assign _cond_data_2188 = (__delay_data_2657__delay_2656__delay_2655_pointer_1562)? 1'sd0 : _cond_data_1311;
  wire signed [16-1:0] _cond_data_2190;
  assign _cond_data_2190 = (__delay_data_2676__delay_2675__delay_2674_pointer_1564)? 1'sd0 : _cond_data_1313;
  wire signed [16-1:0] _cond_data_2192;
  assign _cond_data_2192 = (__delay_data_2693__delay_2692__delay_2691_pointer_1566)? 1'sd0 : _cond_data_1315;
  wire signed [16-1:0] _cond_data_2194;
  assign _cond_data_2194 = (__delay_data_2710__delay_2709__delay_2708_pointer_1568)? 1'sd0 : _cond_data_1317;
  wire signed [16-1:0] _cond_data_2196;
  assign _cond_data_2196 = (__delay_data_2727__delay_2726__delay_2725_pointer_1570)? 1'sd0 : _cond_data_1319;
  wire signed [16-1:0] _cond_data_2198;
  assign _cond_data_2198 = (__delay_data_2744__delay_2743__delay_2742_pointer_1572)? 1'sd0 : _cond_data_1321;
  wire signed [16-1:0] _cond_data_2200;
  assign _cond_data_2200 = (__delay_data_2761__delay_2760__delay_2759_pointer_1574)? 1'sd0 : _cond_data_1323;
  wire signed [16-1:0] _cond_data_2202;
  assign _cond_data_2202 = (__delay_data_2778__delay_2777__delay_2776_pointer_1576)? 1'sd0 : _cond_data_1325;
  wire signed [16-1:0] _cond_data_2204;
  assign _cond_data_2204 = (__delay_data_2795__delay_2794__delay_2793_pointer_1578)? 1'sd0 : _cond_data_1327;
  reg signed [16-1:0] __variable_wdata_743;
  assign mul_35_x_data = __variable_wdata_743;
  reg signed [16-1:0] __variable_wdata_744;
  assign mul_35_y_data = __variable_wdata_744;
  reg [5-1:0] __variable_wdata_745;
  assign mul_35_rshift_data = __variable_wdata_745;
  assign _mul_35_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_35_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_35_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_764;
  assign mul_36_x_data = __variable_wdata_764;
  reg signed [16-1:0] __variable_wdata_765;
  assign mul_36_y_data = __variable_wdata_765;
  reg [5-1:0] __variable_wdata_766;
  assign mul_36_rshift_data = __variable_wdata_766;
  assign _mul_36_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_36_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_36_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_785;
  assign mul_37_x_data = __variable_wdata_785;
  reg signed [16-1:0] __variable_wdata_786;
  assign mul_37_y_data = __variable_wdata_786;
  reg [5-1:0] __variable_wdata_787;
  assign mul_37_rshift_data = __variable_wdata_787;
  assign _mul_37_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_37_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_37_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_806;
  assign mul_38_x_data = __variable_wdata_806;
  reg signed [16-1:0] __variable_wdata_807;
  assign mul_38_y_data = __variable_wdata_807;
  reg [5-1:0] __variable_wdata_808;
  assign mul_38_rshift_data = __variable_wdata_808;
  assign _mul_38_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_38_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_38_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_827;
  assign mul_39_x_data = __variable_wdata_827;
  reg signed [16-1:0] __variable_wdata_828;
  assign mul_39_y_data = __variable_wdata_828;
  reg [5-1:0] __variable_wdata_829;
  assign mul_39_rshift_data = __variable_wdata_829;
  assign _mul_39_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_39_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_39_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_848;
  assign mul_40_x_data = __variable_wdata_848;
  reg signed [16-1:0] __variable_wdata_849;
  assign mul_40_y_data = __variable_wdata_849;
  reg [5-1:0] __variable_wdata_850;
  assign mul_40_rshift_data = __variable_wdata_850;
  assign _mul_40_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_40_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_40_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_869;
  assign mul_41_x_data = __variable_wdata_869;
  reg signed [16-1:0] __variable_wdata_870;
  assign mul_41_y_data = __variable_wdata_870;
  reg [5-1:0] __variable_wdata_871;
  assign mul_41_rshift_data = __variable_wdata_871;
  assign _mul_41_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_41_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_41_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_890;
  assign mul_42_x_data = __variable_wdata_890;
  reg signed [16-1:0] __variable_wdata_891;
  assign mul_42_y_data = __variable_wdata_891;
  reg [5-1:0] __variable_wdata_892;
  assign mul_42_rshift_data = __variable_wdata_892;
  assign _mul_42_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_42_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_42_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_911;
  assign mul_43_x_data = __variable_wdata_911;
  reg signed [16-1:0] __variable_wdata_912;
  assign mul_43_y_data = __variable_wdata_912;
  reg [5-1:0] __variable_wdata_913;
  assign mul_43_rshift_data = __variable_wdata_913;
  assign _mul_43_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_43_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_43_stream_internal_oready;
  reg [1-1:0] __delay_data_2811__delay_2810__delay_2809____variable_951;
  reg [16-1:0] __delay_data_2826__delay_2825__delay_2824_plus_1972;
  reg [6-1:0] __delay_data_2842__delay_2841__delay_2840____variable_946;
  reg [16-1:0] __delay_data_2947__delay_2946__delay_2945_plus_2390;
  reg signed [16-1:0] __delay_data_2963__delay_2962__delay_2961__delay_2960_cond_978;
  reg signed [16-1:0] __delay_data_2985__delay_2984__delay_2983__delay_2982_cond_990;
  reg [16-1:0] __delay_data_3007__delay_3006__delay_3005_plus_2409;
  reg signed [16-1:0] __delay_data_3031__delay_3030__delay_3029__delay_3028_cond_977;
  reg signed [16-1:0] __delay_data_3053__delay_3052__delay_3051__delay_3050_cond_989;
  reg [16-1:0] __delay_data_3075__delay_3074__delay_3073_plus_1991;
  reg [1-1:0] __delay_data_2812__delay_2811__delay_2810____variable_951;
  reg [16-1:0] __delay_data_2827__delay_2826__delay_2825___plus_1972;
  reg [6-1:0] __delay_data_2843__delay_2842__delay_2841____variable_946;
  reg [16-1:0] __delay_data_2948__delay_2947__delay_2946___plus_2390;
  reg signed [16-1:0] __delay_data_2964__delay_2963__delay_2962__delay_2961___cond_978;
  reg signed [16-1:0] __delay_data_2986__delay_2985__delay_2984__delay_2983___cond_990;
  reg [16-1:0] __delay_data_3008__delay_3007__delay_3006___plus_2409;
  reg signed [16-1:0] __delay_data_3032__delay_3031__delay_3030__delay_3029___cond_977;
  reg signed [16-1:0] __delay_data_3054__delay_3053__delay_3052__delay_3051___cond_989;
  reg [16-1:0] __delay_data_3076__delay_3075__delay_3074___plus_1991;
  reg [1-1:0] __delay_data_2813__delay_2812__delay_2811____variable_951;
  reg [16-1:0] __delay_data_2828__delay_2827__delay_2826___plus_1972;
  reg [6-1:0] __delay_data_2844__delay_2843__delay_2842____variable_946;
  reg [16-1:0] __delay_data_2949__delay_2948__delay_2947___plus_2390;
  reg signed [16-1:0] __delay_data_2965__delay_2964__delay_2963__delay_2962___cond_978;
  reg signed [16-1:0] __delay_data_2987__delay_2986__delay_2985__delay_2984___cond_990;
  reg [16-1:0] __delay_data_3009__delay_3008__delay_3007___plus_2409;
  reg signed [16-1:0] __delay_data_3033__delay_3032__delay_3031__delay_3030___cond_977;
  reg signed [16-1:0] __delay_data_3055__delay_3054__delay_3053__delay_3052___cond_989;
  reg [16-1:0] __delay_data_3077__delay_3076__delay_3075___plus_1991;
  reg [1-1:0] __delay_data_2814__delay_2813__delay_2812____variable_951;
  reg [16-1:0] __delay_data_2829__delay_2828__delay_2827___plus_1972;
  reg [6-1:0] __delay_data_2845__delay_2844__delay_2843____variable_946;
  reg [16-1:0] __delay_data_2950__delay_2949__delay_2948___plus_2390;
  reg signed [16-1:0] __delay_data_2966__delay_2965__delay_2964__delay_2963___cond_978;
  reg signed [16-1:0] __delay_data_2988__delay_2987__delay_2986__delay_2985___cond_990;
  reg [16-1:0] __delay_data_3010__delay_3009__delay_3008___plus_2409;
  reg signed [16-1:0] __delay_data_3034__delay_3033__delay_3032__delay_3031___cond_977;
  reg signed [16-1:0] __delay_data_3056__delay_3055__delay_3054__delay_3053___cond_989;
  reg [16-1:0] __delay_data_3078__delay_3077__delay_3076___plus_1991;
  reg [1-1:0] __delay_data_2815__delay_2814__delay_2813____variable_951;
  reg [16-1:0] __delay_data_2830__delay_2829__delay_2828___plus_1972;
  reg [6-1:0] __delay_data_2846__delay_2845__delay_2844____variable_946;
  reg [16-1:0] __delay_data_2951__delay_2950__delay_2949___plus_2390;
  reg signed [16-1:0] __delay_data_2967__delay_2966__delay_2965__delay_2964___cond_978;
  reg signed [16-1:0] __delay_data_2989__delay_2988__delay_2987__delay_2986___cond_990;
  reg [16-1:0] __delay_data_3011__delay_3010__delay_3009___plus_2409;
  reg signed [16-1:0] __delay_data_3035__delay_3034__delay_3033__delay_3032___cond_977;
  reg signed [16-1:0] __delay_data_3057__delay_3056__delay_3055__delay_3054___cond_989;
  reg [16-1:0] __delay_data_3079__delay_3078__delay_3077___plus_1991;
  reg [1-1:0] __delay_data_2816__delay_2815__delay_2814____variable_951;
  reg [16-1:0] __delay_data_2831__delay_2830__delay_2829___plus_1972;
  reg [6-1:0] __delay_data_2847__delay_2846__delay_2845____variable_946;
  reg [16-1:0] __delay_data_2952__delay_2951__delay_2950___plus_2390;
  reg signed [16-1:0] __delay_data_2968__delay_2967__delay_2966__delay_2965___cond_978;
  reg signed [16-1:0] __delay_data_2990__delay_2989__delay_2988__delay_2987___cond_990;
  reg [16-1:0] __delay_data_3012__delay_3011__delay_3010___plus_2409;
  reg signed [16-1:0] __delay_data_3036__delay_3035__delay_3034__delay_3033___cond_977;
  reg signed [16-1:0] __delay_data_3058__delay_3057__delay_3056__delay_3055___cond_989;
  reg [16-1:0] __delay_data_3080__delay_3079__delay_3078___plus_1991;
  reg [1-1:0] __delay_data_2817__delay_2816__delay_2815____variable_951;
  reg [16-1:0] __delay_data_2832__delay_2831__delay_2830___plus_1972;
  reg [6-1:0] __delay_data_2848__delay_2847__delay_2846____variable_946;
  reg [16-1:0] __delay_data_2953__delay_2952__delay_2951___plus_2390;
  reg signed [16-1:0] __delay_data_2969__delay_2968__delay_2967__delay_2966___cond_978;
  reg signed [16-1:0] __delay_data_2991__delay_2990__delay_2989__delay_2988___cond_990;
  reg [16-1:0] __delay_data_3013__delay_3012__delay_3011___plus_2409;
  reg signed [16-1:0] __delay_data_3037__delay_3036__delay_3035__delay_3034___cond_977;
  reg signed [16-1:0] __delay_data_3059__delay_3058__delay_3057__delay_3056___cond_989;
  reg [16-1:0] __delay_data_3081__delay_3080__delay_3079___plus_1991;
  reg [1-1:0] __delay_data_2818__delay_2817__delay_2816____variable_951;
  reg [16-1:0] __delay_data_2833__delay_2832__delay_2831___plus_1972;
  reg [6-1:0] __delay_data_2849__delay_2848__delay_2847____variable_946;
  reg [16-1:0] __delay_data_2954__delay_2953__delay_2952___plus_2390;
  reg signed [16-1:0] __delay_data_2970__delay_2969__delay_2968__delay_2967___cond_978;
  reg signed [16-1:0] __delay_data_2992__delay_2991__delay_2990__delay_2989___cond_990;
  reg [16-1:0] __delay_data_3014__delay_3013__delay_3012___plus_2409;
  reg signed [16-1:0] __delay_data_3038__delay_3037__delay_3036__delay_3035___cond_977;
  reg signed [16-1:0] __delay_data_3060__delay_3059__delay_3058__delay_3057___cond_989;
  reg [16-1:0] __delay_data_3082__delay_3081__delay_3080___plus_1991;
  reg [1-1:0] __delay_data_2819__delay_2818__delay_2817____variable_951;
  reg [16-1:0] __delay_data_2834__delay_2833__delay_2832___plus_1972;
  reg [6-1:0] __delay_data_2850__delay_2849__delay_2848____variable_946;
  reg [16-1:0] __delay_data_2955__delay_2954__delay_2953___plus_2390;
  reg signed [16-1:0] __delay_data_2971__delay_2970__delay_2969__delay_2968___cond_978;
  reg signed [16-1:0] __delay_data_2993__delay_2992__delay_2991__delay_2990___cond_990;
  reg [16-1:0] __delay_data_3015__delay_3014__delay_3013___plus_2409;
  reg signed [16-1:0] __delay_data_3039__delay_3038__delay_3037__delay_3036___cond_977;
  reg signed [16-1:0] __delay_data_3061__delay_3060__delay_3059__delay_3058___cond_989;
  reg [16-1:0] __delay_data_3083__delay_3082__delay_3081___plus_1991;
  wire signed [32-1:0] __substreamoutput_data_1616;
  assign __substreamoutput_data_1616 = mul_8_z_data;
  wire signed [32-1:0] __substreamoutput_data_1635;
  assign __substreamoutput_data_1635 = mul_9_z_data;
  wire signed [32-1:0] __substreamoutput_data_1654;
  assign __substreamoutput_data_1654 = mul_10_z_data;
  wire signed [32-1:0] __substreamoutput_data_1673;
  assign __substreamoutput_data_1673 = mul_11_z_data;
  wire signed [32-1:0] __substreamoutput_data_1692;
  assign __substreamoutput_data_1692 = mul_12_z_data;
  wire signed [32-1:0] __substreamoutput_data_1711;
  assign __substreamoutput_data_1711 = mul_13_z_data;
  wire signed [32-1:0] __substreamoutput_data_1730;
  assign __substreamoutput_data_1730 = mul_14_z_data;
  wire signed [32-1:0] __substreamoutput_data_1749;
  assign __substreamoutput_data_1749 = mul_15_z_data;
  wire signed [32-1:0] __substreamoutput_data_1768;
  assign __substreamoutput_data_1768 = mul_16_z_data;
  wire signed [32-1:0] __substreamoutput_data_1805;
  assign __substreamoutput_data_1805 = mul_17_z_data;
  wire signed [32-1:0] __substreamoutput_data_1824;
  assign __substreamoutput_data_1824 = mul_18_z_data;
  wire signed [32-1:0] __substreamoutput_data_1843;
  assign __substreamoutput_data_1843 = mul_19_z_data;
  wire signed [32-1:0] __substreamoutput_data_1862;
  assign __substreamoutput_data_1862 = mul_20_z_data;
  wire signed [32-1:0] __substreamoutput_data_1881;
  assign __substreamoutput_data_1881 = mul_21_z_data;
  wire signed [32-1:0] __substreamoutput_data_1900;
  assign __substreamoutput_data_1900 = mul_22_z_data;
  wire signed [32-1:0] __substreamoutput_data_1919;
  assign __substreamoutput_data_1919 = mul_23_z_data;
  wire signed [32-1:0] __substreamoutput_data_1938;
  assign __substreamoutput_data_1938 = mul_24_z_data;
  wire signed [32-1:0] __substreamoutput_data_1957;
  assign __substreamoutput_data_1957 = mul_25_z_data;
  reg signed [64-1:0] __variable_wdata_52;
  assign add_tree_4_var0_data = __variable_wdata_52;
  reg signed [64-1:0] __variable_wdata_53;
  assign add_tree_4_var1_data = __variable_wdata_53;
  reg signed [64-1:0] __variable_wdata_54;
  assign add_tree_4_var2_data = __variable_wdata_54;
  reg signed [64-1:0] __variable_wdata_55;
  assign add_tree_4_var3_data = __variable_wdata_55;
  reg signed [64-1:0] __variable_wdata_56;
  assign add_tree_4_var4_data = __variable_wdata_56;
  reg signed [64-1:0] __variable_wdata_57;
  assign add_tree_4_var5_data = __variable_wdata_57;
  reg signed [64-1:0] __variable_wdata_58;
  assign add_tree_4_var6_data = __variable_wdata_58;
  reg signed [64-1:0] __variable_wdata_59;
  assign add_tree_4_var7_data = __variable_wdata_59;
  reg signed [64-1:0] __variable_wdata_60;
  assign add_tree_4_var8_data = __variable_wdata_60;
  reg signed [64-1:0] __variable_wdata_61;
  assign add_tree_4_var9_data = __variable_wdata_61;
  reg signed [64-1:0] __variable_wdata_62;
  assign add_tree_4_var10_data = __variable_wdata_62;
  reg signed [64-1:0] __variable_wdata_63;
  assign add_tree_4_var11_data = __variable_wdata_63;
  reg signed [64-1:0] __variable_wdata_64;
  assign add_tree_4_var12_data = __variable_wdata_64;
  reg signed [64-1:0] __variable_wdata_65;
  assign add_tree_4_var13_data = __variable_wdata_65;
  reg signed [64-1:0] __variable_wdata_66;
  assign add_tree_4_var14_data = __variable_wdata_66;
  reg signed [64-1:0] __variable_wdata_67;
  assign add_tree_4_var15_data = __variable_wdata_67;
  reg signed [64-1:0] __variable_wdata_68;
  assign add_tree_4_var16_data = __variable_wdata_68;
  reg signed [64-1:0] __variable_wdata_69;
  assign add_tree_4_var17_data = __variable_wdata_69;
  assign _add_tree_4_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _add_tree_4_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _add_tree_4_stream_internal_oready;
  wire signed [32-1:0] __substreamoutput_data_2034;
  assign __substreamoutput_data_2034 = mul_26_z_data;
  wire signed [32-1:0] __substreamoutput_data_2053;
  assign __substreamoutput_data_2053 = mul_27_z_data;
  wire signed [32-1:0] __substreamoutput_data_2072;
  assign __substreamoutput_data_2072 = mul_28_z_data;
  wire signed [32-1:0] __substreamoutput_data_2091;
  assign __substreamoutput_data_2091 = mul_29_z_data;
  wire signed [32-1:0] __substreamoutput_data_2110;
  assign __substreamoutput_data_2110 = mul_30_z_data;
  wire signed [32-1:0] __substreamoutput_data_2129;
  assign __substreamoutput_data_2129 = mul_31_z_data;
  wire signed [32-1:0] __substreamoutput_data_2148;
  assign __substreamoutput_data_2148 = mul_32_z_data;
  wire signed [32-1:0] __substreamoutput_data_2167;
  assign __substreamoutput_data_2167 = mul_33_z_data;
  wire signed [32-1:0] __substreamoutput_data_2186;
  assign __substreamoutput_data_2186 = mul_34_z_data;
  wire signed [32-1:0] __substreamoutput_data_2223;
  assign __substreamoutput_data_2223 = mul_35_z_data;
  wire signed [32-1:0] __substreamoutput_data_2242;
  assign __substreamoutput_data_2242 = mul_36_z_data;
  wire signed [32-1:0] __substreamoutput_data_2261;
  assign __substreamoutput_data_2261 = mul_37_z_data;
  wire signed [32-1:0] __substreamoutput_data_2280;
  assign __substreamoutput_data_2280 = mul_38_z_data;
  wire signed [32-1:0] __substreamoutput_data_2299;
  assign __substreamoutput_data_2299 = mul_39_z_data;
  wire signed [32-1:0] __substreamoutput_data_2318;
  assign __substreamoutput_data_2318 = mul_40_z_data;
  wire signed [32-1:0] __substreamoutput_data_2337;
  assign __substreamoutput_data_2337 = mul_41_z_data;
  wire signed [32-1:0] __substreamoutput_data_2356;
  assign __substreamoutput_data_2356 = mul_42_z_data;
  wire signed [32-1:0] __substreamoutput_data_2375;
  assign __substreamoutput_data_2375 = mul_43_z_data;
  reg signed [64-1:0] __variable_wdata_80;
  assign add_tree_5_var0_data = __variable_wdata_80;
  reg signed [64-1:0] __variable_wdata_81;
  assign add_tree_5_var1_data = __variable_wdata_81;
  reg signed [64-1:0] __variable_wdata_82;
  assign add_tree_5_var2_data = __variable_wdata_82;
  reg signed [64-1:0] __variable_wdata_83;
  assign add_tree_5_var3_data = __variable_wdata_83;
  reg signed [64-1:0] __variable_wdata_84;
  assign add_tree_5_var4_data = __variable_wdata_84;
  reg signed [64-1:0] __variable_wdata_85;
  assign add_tree_5_var5_data = __variable_wdata_85;
  reg signed [64-1:0] __variable_wdata_86;
  assign add_tree_5_var6_data = __variable_wdata_86;
  reg signed [64-1:0] __variable_wdata_87;
  assign add_tree_5_var7_data = __variable_wdata_87;
  reg signed [64-1:0] __variable_wdata_88;
  assign add_tree_5_var8_data = __variable_wdata_88;
  reg signed [64-1:0] __variable_wdata_89;
  assign add_tree_5_var9_data = __variable_wdata_89;
  reg signed [64-1:0] __variable_wdata_90;
  assign add_tree_5_var10_data = __variable_wdata_90;
  reg signed [64-1:0] __variable_wdata_91;
  assign add_tree_5_var11_data = __variable_wdata_91;
  reg signed [64-1:0] __variable_wdata_92;
  assign add_tree_5_var12_data = __variable_wdata_92;
  reg signed [64-1:0] __variable_wdata_93;
  assign add_tree_5_var13_data = __variable_wdata_93;
  reg signed [64-1:0] __variable_wdata_94;
  assign add_tree_5_var14_data = __variable_wdata_94;
  reg signed [64-1:0] __variable_wdata_95;
  assign add_tree_5_var15_data = __variable_wdata_95;
  reg signed [64-1:0] __variable_wdata_96;
  assign add_tree_5_var16_data = __variable_wdata_96;
  reg signed [64-1:0] __variable_wdata_97;
  assign add_tree_5_var17_data = __variable_wdata_97;
  assign _add_tree_5_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _add_tree_5_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _add_tree_5_stream_internal_oready;
  reg [1-1:0] __delay_data_2820__delay_2819__delay_2818____variable_951;
  reg [16-1:0] __delay_data_2835__delay_2834__delay_2833___plus_1972;
  reg [6-1:0] __delay_data_2851__delay_2850__delay_2849____variable_946;
  reg [16-1:0] __delay_data_2956__delay_2955__delay_2954___plus_2390;
  reg signed [16-1:0] __delay_data_2972__delay_2971__delay_2970__delay_2969___cond_978;
  reg signed [16-1:0] __delay_data_2994__delay_2993__delay_2992__delay_2991___cond_990;
  reg [16-1:0] __delay_data_3016__delay_3015__delay_3014___plus_2409;
  reg signed [16-1:0] __delay_data_3040__delay_3039__delay_3038__delay_3037___cond_977;
  reg signed [16-1:0] __delay_data_3062__delay_3061__delay_3060__delay_3059___cond_989;
  reg [16-1:0] __delay_data_3084__delay_3083__delay_3082___plus_1991;
  reg [1-1:0] __delay_data_2821__delay_2820__delay_2819____variable_951;
  reg [16-1:0] __delay_data_2836__delay_2835__delay_2834___plus_1972;
  reg [6-1:0] __delay_data_2852__delay_2851__delay_2850____variable_946;
  reg [16-1:0] __delay_data_2957__delay_2956__delay_2955___plus_2390;
  reg signed [16-1:0] __delay_data_2973__delay_2972__delay_2971__delay_2970___cond_978;
  reg signed [16-1:0] __delay_data_2995__delay_2994__delay_2993__delay_2992___cond_990;
  reg [16-1:0] __delay_data_3017__delay_3016__delay_3015___plus_2409;
  reg signed [16-1:0] __delay_data_3041__delay_3040__delay_3039__delay_3038___cond_977;
  reg signed [16-1:0] __delay_data_3063__delay_3062__delay_3061__delay_3060___cond_989;
  reg [16-1:0] __delay_data_3085__delay_3084__delay_3083___plus_1991;
  reg [1-1:0] __delay_data_2822__delay_2821__delay_2820____variable_951;
  reg [16-1:0] __delay_data_2837__delay_2836__delay_2835___plus_1972;
  reg [6-1:0] __delay_data_2853__delay_2852__delay_2851____variable_946;
  reg [16-1:0] __delay_data_2958__delay_2957__delay_2956___plus_2390;
  reg signed [16-1:0] __delay_data_2974__delay_2973__delay_2972__delay_2971___cond_978;
  reg signed [16-1:0] __delay_data_2996__delay_2995__delay_2994__delay_2993___cond_990;
  reg [16-1:0] __delay_data_3018__delay_3017__delay_3016___plus_2409;
  reg signed [16-1:0] __delay_data_3042__delay_3041__delay_3040__delay_3039___cond_977;
  reg signed [16-1:0] __delay_data_3064__delay_3063__delay_3062__delay_3061___cond_989;
  reg [16-1:0] __delay_data_3086__delay_3085__delay_3084___plus_1991;
  reg [1-1:0] __delay_data_2823__delay_2822__delay_2821____variable_951;
  reg [16-1:0] __delay_data_2838__delay_2837__delay_2836___plus_1972;
  reg [6-1:0] __delay_data_2854__delay_2853__delay_2852____variable_946;
  reg [16-1:0] __delay_data_2959__delay_2958__delay_2957___plus_2390;
  reg signed [16-1:0] __delay_data_2975__delay_2974__delay_2973__delay_2972___cond_978;
  reg signed [16-1:0] __delay_data_2997__delay_2996__delay_2995__delay_2994___cond_990;
  reg [16-1:0] __delay_data_3019__delay_3018__delay_3017___plus_2409;
  reg signed [16-1:0] __delay_data_3043__delay_3042__delay_3041__delay_3040___cond_977;
  reg signed [16-1:0] __delay_data_3065__delay_3064__delay_3063__delay_3062___cond_989;
  reg [16-1:0] __delay_data_3087__delay_3086__delay_3085___plus_1991;
  wire signed [64-1:0] __substreamoutput_data_1959;
  assign __substreamoutput_data_1959 = add_tree_4_sum_data;
  reg [1-1:0] __variable_wdata_15;
  assign acc_0__reduce_reset_data = __variable_wdata_15;
  reg signed [64-1:0] __variable_wdata_0;
  assign acc_0_x_data = __variable_wdata_0;
  reg [7-1:0] __variable_wdata_1;
  assign acc_0_rshift_data = __variable_wdata_1;
  reg [32-1:0] __variable_wdata_2;
  assign acc_0_size_data = __variable_wdata_2;
  wire signed [64-1:0] __substreamoutput_data_2377;
  assign __substreamoutput_data_2377 = add_tree_5_sum_data;
  reg [1-1:0] __variable_wdata_37;
  assign acc_1__reduce_reset_data = __variable_wdata_37;
  reg signed [64-1:0] __variable_wdata_22;
  assign acc_1_x_data = __variable_wdata_22;
  reg [7-1:0] __variable_wdata_23;
  assign acc_1_rshift_data = __variable_wdata_23;
  reg [32-1:0] __variable_wdata_24;
  assign acc_1_size_data = __variable_wdata_24;
  reg signed [16-1:0] __delay_data_2976__delay_2975__delay_2974__delay_2973___cond_978;
  reg signed [16-1:0] __delay_data_2998__delay_2997__delay_2996__delay_2995___cond_990;
  reg [16-1:0] __delay_data_3020__delay_3019__delay_3018___plus_2409;
  reg signed [16-1:0] __delay_data_3044__delay_3043__delay_3042__delay_3041___cond_977;
  reg signed [16-1:0] __delay_data_3066__delay_3065__delay_3064__delay_3063___cond_989;
  reg [16-1:0] __delay_data_3088__delay_3087__delay_3086___plus_1991;
  reg signed [16-1:0] __delay_data_2977__delay_2976__delay_2975__delay_2974___cond_978;
  reg signed [16-1:0] __delay_data_2999__delay_2998__delay_2997__delay_2996___cond_990;
  reg [16-1:0] __delay_data_3021__delay_3020__delay_3019___plus_2409;
  reg signed [16-1:0] __delay_data_3045__delay_3044__delay_3043__delay_3042___cond_977;
  reg signed [16-1:0] __delay_data_3067__delay_3066__delay_3065__delay_3064___cond_989;
  reg [16-1:0] __delay_data_3089__delay_3088__delay_3087___plus_1991;
  reg signed [16-1:0] __delay_data_2978__delay_2977__delay_2976__delay_2975___cond_978;
  reg signed [16-1:0] __delay_data_3000__delay_2999__delay_2998__delay_2997___cond_990;
  reg [16-1:0] __delay_data_3022__delay_3021__delay_3020___plus_2409;
  reg signed [16-1:0] __delay_data_3046__delay_3045__delay_3044__delay_3043___cond_977;
  reg signed [16-1:0] __delay_data_3068__delay_3067__delay_3066__delay_3065___cond_989;
  reg [16-1:0] __delay_data_3090__delay_3089__delay_3088___plus_1991;
  reg signed [16-1:0] __delay_data_2979__delay_2978__delay_2977__delay_2976___cond_978;
  reg signed [16-1:0] __delay_data_3001__delay_3000__delay_2999__delay_2998___cond_990;
  reg [16-1:0] __delay_data_3023__delay_3022__delay_3021___plus_2409;
  reg signed [16-1:0] __delay_data_3047__delay_3046__delay_3045__delay_3044___cond_977;
  reg signed [16-1:0] __delay_data_3069__delay_3068__delay_3067__delay_3066___cond_989;
  reg [16-1:0] __delay_data_3091__delay_3090__delay_3089___plus_1991;
  reg signed [16-1:0] __delay_data_2980__delay_2979__delay_2978__delay_2977___cond_978;
  reg signed [16-1:0] __delay_data_3002__delay_3001__delay_3000__delay_2999___cond_990;
  reg [16-1:0] __delay_data_3024__delay_3023__delay_3022___plus_2409;
  reg signed [16-1:0] __delay_data_3048__delay_3047__delay_3046__delay_3045___cond_977;
  reg signed [16-1:0] __delay_data_3070__delay_3069__delay_3068__delay_3067___cond_989;
  reg [16-1:0] __delay_data_3092__delay_3091__delay_3090___plus_1991;
  reg signed [16-1:0] __delay_data_2981__delay_2980__delay_2979__delay_2978___cond_978;
  reg signed [16-1:0] __delay_data_3003__delay_3002__delay_3001__delay_3000___cond_990;
  reg [16-1:0] __delay_data_3025__delay_3024__delay_3023___plus_2409;
  reg signed [16-1:0] __delay_data_3049__delay_3048__delay_3047__delay_3046___cond_977;
  reg signed [16-1:0] __delay_data_3071__delay_3070__delay_3069__delay_3068___cond_989;
  reg [16-1:0] __delay_data_3093__delay_3092__delay_3091___plus_1991;
  wire signed [64-1:0] __substreamoutput_data_1973;
  assign __substreamoutput_data_1973 = acc_0_sum_data;
  wire [1-1:0] __substreamoutput_data_1974;
  assign __substreamoutput_data_1974 = acc_0_valid_data;
  reg signed [64-1:0] _plus_data_1975;
  wire signed [64-1:0] __substreamoutput_data_2391;
  assign __substreamoutput_data_2391 = acc_1_sum_data;
  reg signed [64-1:0] _plus_data_2393;
  reg signed [16-1:0] __delay_data_3004__delay_3003__delay_3002__delay_3001___cond_990;
  reg [16-1:0] __delay_data_3026__delay_3025__delay_3024___plus_2409;
  reg signed [16-1:0] __delay_data_3072__delay_3071__delay_3070__delay_3069___cond_989;
  reg [16-1:0] __delay_data_3094__delay_3093__delay_3092___plus_1991;
  reg [1-1:0] __delay_data_3096__substreamoutput_1974;
  reg signed [64-1:0] __variable_wdata_108;
  assign mul_rshift_round_clip_6_x_data = __variable_wdata_108;
  reg signed [16-1:0] __variable_wdata_109;
  assign mul_rshift_round_clip_6_y_data = __variable_wdata_109;
  reg [7-1:0] __variable_wdata_110;
  assign mul_rshift_round_clip_6_rshift_data = __variable_wdata_110;
  reg signed [64-1:0] __variable_wdata_142;
  assign mul_rshift_round_clip_7_x_data = __variable_wdata_142;
  reg signed [16-1:0] __variable_wdata_143;
  assign mul_rshift_round_clip_7_y_data = __variable_wdata_143;
  reg [7-1:0] __variable_wdata_144;
  assign mul_rshift_round_clip_7_rshift_data = __variable_wdata_144;
  assign _stream_conv2d_4_stream_internal_oready = ((_stream_conv2d_4_busy)? _mul_rshift_round_clip_7_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_rshift_round_clip_6_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _acc_1_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _acc_0_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _add_tree_5_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _add_tree_4_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_43_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_42_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_41_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_40_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_39_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_38_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_37_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_36_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_35_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_34_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_33_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_32_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_31_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_30_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_29_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_28_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_27_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_26_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_25_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_24_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_23_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_22_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_21_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_20_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_19_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_18_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_17_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_16_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_15_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_14_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_13_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_12_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_11_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_10_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_9_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_8_stream_internal_oready : 1) && 1)))))))))))))))))))))))))))))))))))))))));
  reg [1-1:0] __delay_data_3097__delay_3096__substreamoutput_1974;
  reg [1-1:0] __delay_data_3098__delay_3097____substreamoutput_1974;
  reg [1-1:0] __delay_data_3099__delay_3098____substreamoutput_1974;
  reg [1-1:0] __delay_data_3100__delay_3099____substreamoutput_1974;
  reg [1-1:0] __delay_data_3101__delay_3100____substreamoutput_1974;
  reg [1-1:0] __delay_data_3102__delay_3101____substreamoutput_1974;
  reg [1-1:0] __delay_data_3103__delay_3102____substreamoutput_1974;
  reg [1-1:0] __delay_data_3104__delay_3103____substreamoutput_1974;
  reg [1-1:0] __delay_data_3105__delay_3104____substreamoutput_1974;
  wire signed [16-1:0] __substreamoutput_data_1992;
  assign __substreamoutput_data_1992 = mul_rshift_round_clip_6_z_data;
  reg [1-1:0] _greaterthan_data_1994;
  wire signed [16-1:0] __substreamoutput_data_2410;
  assign __substreamoutput_data_2410 = mul_rshift_round_clip_7_z_data;
  reg [1-1:0] _greaterthan_data_2412;
  reg signed [16-1:0] __delay_data_3027__substreamoutput_2410;
  reg signed [16-1:0] __delay_data_3095__substreamoutput_1992;
  reg [1-1:0] __delay_data_3106__delay_3105____substreamoutput_1974;
  reg signed [16-1:0] _cond_data_1996;
  reg signed [16-1:0] _cond_data_2414;
  reg [1-1:0] __delay_data_3107__delay_3106____substreamoutput_1974;
  wire signed [16-1:0] _reinterpretcast_src_1997;
  assign _reinterpretcast_src_1997 = _cond_data_1996;
  wire signed [16-1:0] _reinterpretcast_data_1997;
  assign _reinterpretcast_data_1997 = _reinterpretcast_src_1997;
  wire signed [16-1:0] _reinterpretcast_src_2415;
  assign _reinterpretcast_src_2415 = _cond_data_2414;
  wire signed [16-1:0] _reinterpretcast_data_2415;
  assign _reinterpretcast_data_2415 = _reinterpretcast_src_2415;
  wire [32-1:0] _cat_data_2416;
  assign _cat_data_2416 = { _reinterpretcast_data_2415, _reinterpretcast_data_1997 };
  wire [32-1:0] stream_conv2d_4_sink_89_data;
  assign stream_conv2d_4_sink_89_data = _cat_data_2416;
  wire [1-1:0] stream_conv2d_4_sink_90_data;
  assign stream_conv2d_4_sink_90_data = __delay_data_3107__delay_3106____substreamoutput_1974;
  wire _set_flag_272;
  assign _set_flag_272 = conv2d_4_comp_fsm == 3;
  reg [6-1:0] __variable_wdata_946;
  assign stream_conv2d_4_parameter_0_data = __variable_wdata_946;
  wire _set_flag_273;
  assign _set_flag_273 = conv2d_4_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_947;
  assign stream_conv2d_4_parameter_1_data = __variable_wdata_947;
  wire _set_flag_274;
  assign _set_flag_274 = conv2d_4_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_948;
  assign stream_conv2d_4_parameter_2_data = __variable_wdata_948;
  wire _set_flag_275;
  assign _set_flag_275 = conv2d_4_comp_fsm == 3;
  reg [9-1:0] __variable_wdata_949;
  assign stream_conv2d_4_parameter_3_data = __variable_wdata_949;
  wire _set_flag_276;
  assign _set_flag_276 = conv2d_4_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_950;
  assign stream_conv2d_4_parameter_4_data = __variable_wdata_950;
  wire _set_flag_277;
  assign _set_flag_277 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_967;
  assign stream_conv2d_4_parameter_6_data = __variable_wdata_967;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_3;
  wire _set_flag_278;
  assign _set_flag_278 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id18_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? _stream_conv2d_4_source_7_source_ram_raddr : 'hx;
  assign ram_w32_l128_id18_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_279 = 1;
  wire [_tmp_279-1:0] _tmp_280;
  assign _tmp_280 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1);
  reg [_tmp_279-1:0] __tmp_280_1;
  assign _stream_conv2d_4_source_7_source_ram_rdata = (_stream_conv2d_4_source_7_source_sel == 1)? ram_w32_l128_id18_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_968;
  assign stream_conv2d_4_source_7_data = __variable_wdata_968;
  reg [32-1:0] _stream_conv2d_4_source_7_source_pat_fsm_0;
  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_7_source_pat_all_offset;
  assign _stream_conv2d_4_source_7_source_pat_all_offset = _stream_conv2d_4_source_7_source_offset_buf + _source_stream_conv2d_4_source_7_pat_cur_offset_0 + _source_stream_conv2d_4_source_7_pat_cur_offset_1 + _source_stream_conv2d_4_source_7_pat_cur_offset_2 + _source_stream_conv2d_4_source_7_pat_cur_offset_3;
  wire _set_flag_281;
  assign _set_flag_281 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_979;
  assign stream_conv2d_4_parameter_8_data = __variable_wdata_979;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_3;
  wire _set_flag_282;
  assign _set_flag_282 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id19_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? _stream_conv2d_4_source_9_source_ram_raddr : 'hx;
  assign ram_w32_l128_id19_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_283 = 1;
  wire [_tmp_283-1:0] _tmp_284;
  assign _tmp_284 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2);
  reg [_tmp_283-1:0] __tmp_284_1;
  assign _stream_conv2d_4_source_9_source_ram_rdata = (_stream_conv2d_4_source_9_source_sel == 2)? ram_w32_l128_id19_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_980;
  assign stream_conv2d_4_source_9_data = __variable_wdata_980;
  reg [32-1:0] _stream_conv2d_4_source_9_source_pat_fsm_1;
  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_9_source_pat_all_offset;
  assign _stream_conv2d_4_source_9_source_pat_all_offset = _stream_conv2d_4_source_9_source_offset_buf + _source_stream_conv2d_4_source_9_pat_cur_offset_0 + _source_stream_conv2d_4_source_9_pat_cur_offset_1 + _source_stream_conv2d_4_source_9_pat_cur_offset_2 + _source_stream_conv2d_4_source_9_pat_cur_offset_3;
  wire _set_flag_285;
  assign _set_flag_285 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_991;
  assign stream_conv2d_4_parameter_10_data = __variable_wdata_991;
  wire _set_flag_286;
  assign _set_flag_286 = conv2d_4_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_992;
  assign stream_conv2d_4_source_11_data = __variable_wdata_992;
  wire _set_flag_287;
  assign _set_flag_287 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1003;
  assign stream_conv2d_4_parameter_12_data = __variable_wdata_1003;
  wire _set_flag_288;
  assign _set_flag_288 = conv2d_4_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_1004;
  assign stream_conv2d_4_source_13_data = __variable_wdata_1004;
  wire _set_flag_289;
  assign _set_flag_289 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1015;
  assign stream_conv2d_4_parameter_14_data = __variable_wdata_1015;
  wire _set_flag_290;
  assign _set_flag_290 = conv2d_4_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_1016;
  assign stream_conv2d_4_source_15_data = __variable_wdata_1016;
  wire _set_flag_291;
  assign _set_flag_291 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1027;
  assign stream_conv2d_4_parameter_16_data = __variable_wdata_1027;
  wire _set_flag_292;
  assign _set_flag_292 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1028;
  assign stream_conv2d_4_parameter_17_data = __variable_wdata_1028;
  wire _set_flag_293;
  assign _set_flag_293 = conv2d_4_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_1029;
  assign stream_conv2d_4_parameter_18_data = __variable_wdata_1029;
  wire _set_flag_294;
  assign _set_flag_294 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1030;
  assign stream_conv2d_4_parameter_19_data = __variable_wdata_1030;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_3;
  wire _set_flag_295;
  assign _set_flag_295 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? _stream_conv2d_4_source_20_source_ram_raddr : 'hx;
  assign ram_w32_l512_id0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_296 = 1;
  wire [_tmp_296-1:0] _tmp_297;
  assign _tmp_297 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3);
  reg [_tmp_296-1:0] __tmp_297_1;
  assign _stream_conv2d_4_source_20_source_ram_rdata = (_stream_conv2d_4_source_20_source_sel == 3)? ram_w32_l512_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1031;
  assign stream_conv2d_4_source_20_data = __variable_wdata_1031;
  reg [32-1:0] _stream_conv2d_4_source_20_source_pat_fsm_2;
  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_20_source_pat_all_offset;
  assign _stream_conv2d_4_source_20_source_pat_all_offset = _stream_conv2d_4_source_20_source_offset_buf + _source_stream_conv2d_4_source_20_pat_cur_offset_0 + _source_stream_conv2d_4_source_20_pat_cur_offset_1 + _source_stream_conv2d_4_source_20_pat_cur_offset_2 + _source_stream_conv2d_4_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_3;
  wire _set_flag_298;
  assign _set_flag_298 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? _stream_conv2d_4_source_21_source_ram_raddr : 'hx;
  assign ram_w32_l512_id1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_299 = 1;
  wire [_tmp_299-1:0] _tmp_300;
  assign _tmp_300 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4);
  reg [_tmp_299-1:0] __tmp_300_1;
  assign _stream_conv2d_4_source_21_source_ram_rdata = (_stream_conv2d_4_source_21_source_sel == 4)? ram_w32_l512_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1032;
  assign stream_conv2d_4_source_21_data = __variable_wdata_1032;
  reg [32-1:0] _stream_conv2d_4_source_21_source_pat_fsm_3;
  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_21_source_pat_all_offset;
  assign _stream_conv2d_4_source_21_source_pat_all_offset = _stream_conv2d_4_source_21_source_offset_buf + _source_stream_conv2d_4_source_21_pat_cur_offset_0 + _source_stream_conv2d_4_source_21_pat_cur_offset_1 + _source_stream_conv2d_4_source_21_pat_cur_offset_2 + _source_stream_conv2d_4_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_3;
  wire _set_flag_301;
  assign _set_flag_301 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id2_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? _stream_conv2d_4_source_22_source_ram_raddr : 'hx;
  assign ram_w32_l512_id2_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_302 = 1;
  wire [_tmp_302-1:0] _tmp_303;
  assign _tmp_303 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5);
  reg [_tmp_302-1:0] __tmp_303_1;
  assign _stream_conv2d_4_source_22_source_ram_rdata = (_stream_conv2d_4_source_22_source_sel == 5)? ram_w32_l512_id2_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1033;
  assign stream_conv2d_4_source_22_data = __variable_wdata_1033;
  reg [32-1:0] _stream_conv2d_4_source_22_source_pat_fsm_4;
  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_22_source_pat_all_offset;
  assign _stream_conv2d_4_source_22_source_pat_all_offset = _stream_conv2d_4_source_22_source_offset_buf + _source_stream_conv2d_4_source_22_pat_cur_offset_0 + _source_stream_conv2d_4_source_22_pat_cur_offset_1 + _source_stream_conv2d_4_source_22_pat_cur_offset_2 + _source_stream_conv2d_4_source_22_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_3;
  wire _set_flag_304;
  assign _set_flag_304 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id3_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? _stream_conv2d_4_source_23_source_ram_raddr : 'hx;
  assign ram_w32_l512_id3_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_305 = 1;
  wire [_tmp_305-1:0] _tmp_306;
  assign _tmp_306 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6);
  reg [_tmp_305-1:0] __tmp_306_1;
  assign _stream_conv2d_4_source_23_source_ram_rdata = (_stream_conv2d_4_source_23_source_sel == 6)? ram_w32_l512_id3_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1034;
  assign stream_conv2d_4_source_23_data = __variable_wdata_1034;
  reg [32-1:0] _stream_conv2d_4_source_23_source_pat_fsm_5;
  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_23_source_pat_all_offset;
  assign _stream_conv2d_4_source_23_source_pat_all_offset = _stream_conv2d_4_source_23_source_offset_buf + _source_stream_conv2d_4_source_23_pat_cur_offset_0 + _source_stream_conv2d_4_source_23_pat_cur_offset_1 + _source_stream_conv2d_4_source_23_pat_cur_offset_2 + _source_stream_conv2d_4_source_23_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_3;
  wire _set_flag_307;
  assign _set_flag_307 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id4_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? _stream_conv2d_4_source_24_source_ram_raddr : 'hx;
  assign ram_w32_l512_id4_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_308 = 1;
  wire [_tmp_308-1:0] _tmp_309;
  assign _tmp_309 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7);
  reg [_tmp_308-1:0] __tmp_309_1;
  assign _stream_conv2d_4_source_24_source_ram_rdata = (_stream_conv2d_4_source_24_source_sel == 7)? ram_w32_l512_id4_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1035;
  assign stream_conv2d_4_source_24_data = __variable_wdata_1035;
  reg [32-1:0] _stream_conv2d_4_source_24_source_pat_fsm_6;
  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_24_source_pat_all_offset;
  assign _stream_conv2d_4_source_24_source_pat_all_offset = _stream_conv2d_4_source_24_source_offset_buf + _source_stream_conv2d_4_source_24_pat_cur_offset_0 + _source_stream_conv2d_4_source_24_pat_cur_offset_1 + _source_stream_conv2d_4_source_24_pat_cur_offset_2 + _source_stream_conv2d_4_source_24_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_3;
  wire _set_flag_310;
  assign _set_flag_310 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id5_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? _stream_conv2d_4_source_25_source_ram_raddr : 'hx;
  assign ram_w32_l512_id5_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_311 = 1;
  wire [_tmp_311-1:0] _tmp_312;
  assign _tmp_312 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8);
  reg [_tmp_311-1:0] __tmp_312_1;
  assign _stream_conv2d_4_source_25_source_ram_rdata = (_stream_conv2d_4_source_25_source_sel == 8)? ram_w32_l512_id5_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1036;
  assign stream_conv2d_4_source_25_data = __variable_wdata_1036;
  reg [32-1:0] _stream_conv2d_4_source_25_source_pat_fsm_7;
  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_25_source_pat_all_offset;
  assign _stream_conv2d_4_source_25_source_pat_all_offset = _stream_conv2d_4_source_25_source_offset_buf + _source_stream_conv2d_4_source_25_pat_cur_offset_0 + _source_stream_conv2d_4_source_25_pat_cur_offset_1 + _source_stream_conv2d_4_source_25_pat_cur_offset_2 + _source_stream_conv2d_4_source_25_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_3;
  wire _set_flag_313;
  assign _set_flag_313 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id6_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? _stream_conv2d_4_source_26_source_ram_raddr : 'hx;
  assign ram_w32_l512_id6_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_314 = 1;
  wire [_tmp_314-1:0] _tmp_315;
  assign _tmp_315 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9);
  reg [_tmp_314-1:0] __tmp_315_1;
  assign _stream_conv2d_4_source_26_source_ram_rdata = (_stream_conv2d_4_source_26_source_sel == 9)? ram_w32_l512_id6_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1037;
  assign stream_conv2d_4_source_26_data = __variable_wdata_1037;
  reg [32-1:0] _stream_conv2d_4_source_26_source_pat_fsm_8;
  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_26_source_pat_all_offset;
  assign _stream_conv2d_4_source_26_source_pat_all_offset = _stream_conv2d_4_source_26_source_offset_buf + _source_stream_conv2d_4_source_26_pat_cur_offset_0 + _source_stream_conv2d_4_source_26_pat_cur_offset_1 + _source_stream_conv2d_4_source_26_pat_cur_offset_2 + _source_stream_conv2d_4_source_26_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_3;
  wire _set_flag_316;
  assign _set_flag_316 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id7_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? _stream_conv2d_4_source_27_source_ram_raddr : 'hx;
  assign ram_w32_l512_id7_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_317 = 1;
  wire [_tmp_317-1:0] _tmp_318;
  assign _tmp_318 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10);
  reg [_tmp_317-1:0] __tmp_318_1;
  assign _stream_conv2d_4_source_27_source_ram_rdata = (_stream_conv2d_4_source_27_source_sel == 10)? ram_w32_l512_id7_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1038;
  assign stream_conv2d_4_source_27_data = __variable_wdata_1038;
  reg [32-1:0] _stream_conv2d_4_source_27_source_pat_fsm_9;
  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_27_source_pat_all_offset;
  assign _stream_conv2d_4_source_27_source_pat_all_offset = _stream_conv2d_4_source_27_source_offset_buf + _source_stream_conv2d_4_source_27_pat_cur_offset_0 + _source_stream_conv2d_4_source_27_pat_cur_offset_1 + _source_stream_conv2d_4_source_27_pat_cur_offset_2 + _source_stream_conv2d_4_source_27_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_3;
  wire _set_flag_319;
  assign _set_flag_319 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l512_id8_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? _stream_conv2d_4_source_28_source_ram_raddr : 'hx;
  assign ram_w32_l512_id8_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_320 = 1;
  wire [_tmp_320-1:0] _tmp_321;
  assign _tmp_321 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11);
  reg [_tmp_320-1:0] __tmp_321_1;
  assign _stream_conv2d_4_source_28_source_ram_rdata = (_stream_conv2d_4_source_28_source_sel == 11)? ram_w32_l512_id8_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1039;
  assign stream_conv2d_4_source_28_data = __variable_wdata_1039;
  reg [32-1:0] _stream_conv2d_4_source_28_source_pat_fsm_10;
  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_28_source_pat_all_offset;
  assign _stream_conv2d_4_source_28_source_pat_all_offset = _stream_conv2d_4_source_28_source_offset_buf + _source_stream_conv2d_4_source_28_pat_cur_offset_0 + _source_stream_conv2d_4_source_28_pat_cur_offset_1 + _source_stream_conv2d_4_source_28_pat_cur_offset_2 + _source_stream_conv2d_4_source_28_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_3;
  wire _set_flag_322;
  assign _set_flag_322 = conv2d_4_comp_fsm == 3;
  localparam _tmp_323 = 1;
  wire [_tmp_323-1:0] _tmp_324;
  assign _tmp_324 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12);
  reg [_tmp_323-1:0] __tmp_324_1;
  assign _stream_conv2d_4_source_29_source_ram_rdata = (_stream_conv2d_4_source_29_source_sel == 12)? ram_w32_l128_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1328;
  assign stream_conv2d_4_source_29_data = __variable_wdata_1328;
  reg [32-1:0] _stream_conv2d_4_source_29_source_pat_fsm_11;
  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_29_source_pat_all_offset;
  assign _stream_conv2d_4_source_29_source_pat_all_offset = _stream_conv2d_4_source_29_source_offset_buf + _source_stream_conv2d_4_source_29_pat_cur_offset_0 + _source_stream_conv2d_4_source_29_pat_cur_offset_1 + _source_stream_conv2d_4_source_29_pat_cur_offset_2 + _source_stream_conv2d_4_source_29_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_3;
  wire _set_flag_325;
  assign _set_flag_325 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? _stream_conv2d_4_source_30_source_ram_raddr : 'hx;
  assign ram_w32_l128_id1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_326 = 1;
  wire [_tmp_326-1:0] _tmp_327;
  assign _tmp_327 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13);
  reg [_tmp_326-1:0] __tmp_327_1;
  assign _stream_conv2d_4_source_30_source_ram_rdata = (_stream_conv2d_4_source_30_source_sel == 13)? ram_w32_l128_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1329;
  assign stream_conv2d_4_source_30_data = __variable_wdata_1329;
  reg [32-1:0] _stream_conv2d_4_source_30_source_pat_fsm_12;
  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_30_source_pat_all_offset;
  assign _stream_conv2d_4_source_30_source_pat_all_offset = _stream_conv2d_4_source_30_source_offset_buf + _source_stream_conv2d_4_source_30_pat_cur_offset_0 + _source_stream_conv2d_4_source_30_pat_cur_offset_1 + _source_stream_conv2d_4_source_30_pat_cur_offset_2 + _source_stream_conv2d_4_source_30_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_3;
  wire _set_flag_328;
  assign _set_flag_328 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id2_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? _stream_conv2d_4_source_31_source_ram_raddr : 'hx;
  assign ram_w32_l128_id2_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_329 = 1;
  wire [_tmp_329-1:0] _tmp_330;
  assign _tmp_330 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14);
  reg [_tmp_329-1:0] __tmp_330_1;
  assign _stream_conv2d_4_source_31_source_ram_rdata = (_stream_conv2d_4_source_31_source_sel == 14)? ram_w32_l128_id2_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1330;
  assign stream_conv2d_4_source_31_data = __variable_wdata_1330;
  reg [32-1:0] _stream_conv2d_4_source_31_source_pat_fsm_13;
  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_31_source_pat_all_offset;
  assign _stream_conv2d_4_source_31_source_pat_all_offset = _stream_conv2d_4_source_31_source_offset_buf + _source_stream_conv2d_4_source_31_pat_cur_offset_0 + _source_stream_conv2d_4_source_31_pat_cur_offset_1 + _source_stream_conv2d_4_source_31_pat_cur_offset_2 + _source_stream_conv2d_4_source_31_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_3;
  wire _set_flag_331;
  assign _set_flag_331 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id3_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? _stream_conv2d_4_source_32_source_ram_raddr : 'hx;
  assign ram_w32_l128_id3_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_332 = 1;
  wire [_tmp_332-1:0] _tmp_333;
  assign _tmp_333 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15);
  reg [_tmp_332-1:0] __tmp_333_1;
  assign _stream_conv2d_4_source_32_source_ram_rdata = (_stream_conv2d_4_source_32_source_sel == 15)? ram_w32_l128_id3_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1331;
  assign stream_conv2d_4_source_32_data = __variable_wdata_1331;
  reg [32-1:0] _stream_conv2d_4_source_32_source_pat_fsm_14;
  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_32_source_pat_all_offset;
  assign _stream_conv2d_4_source_32_source_pat_all_offset = _stream_conv2d_4_source_32_source_offset_buf + _source_stream_conv2d_4_source_32_pat_cur_offset_0 + _source_stream_conv2d_4_source_32_pat_cur_offset_1 + _source_stream_conv2d_4_source_32_pat_cur_offset_2 + _source_stream_conv2d_4_source_32_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_3;
  wire _set_flag_334;
  assign _set_flag_334 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id4_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? _stream_conv2d_4_source_33_source_ram_raddr : 'hx;
  assign ram_w32_l128_id4_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_335 = 1;
  wire [_tmp_335-1:0] _tmp_336;
  assign _tmp_336 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16);
  reg [_tmp_335-1:0] __tmp_336_1;
  assign _stream_conv2d_4_source_33_source_ram_rdata = (_stream_conv2d_4_source_33_source_sel == 16)? ram_w32_l128_id4_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1332;
  assign stream_conv2d_4_source_33_data = __variable_wdata_1332;
  reg [32-1:0] _stream_conv2d_4_source_33_source_pat_fsm_15;
  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_33_source_pat_all_offset;
  assign _stream_conv2d_4_source_33_source_pat_all_offset = _stream_conv2d_4_source_33_source_offset_buf + _source_stream_conv2d_4_source_33_pat_cur_offset_0 + _source_stream_conv2d_4_source_33_pat_cur_offset_1 + _source_stream_conv2d_4_source_33_pat_cur_offset_2 + _source_stream_conv2d_4_source_33_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_3;
  wire _set_flag_337;
  assign _set_flag_337 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id5_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? _stream_conv2d_4_source_34_source_ram_raddr : 'hx;
  assign ram_w32_l128_id5_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_338 = 1;
  wire [_tmp_338-1:0] _tmp_339;
  assign _tmp_339 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17);
  reg [_tmp_338-1:0] __tmp_339_1;
  assign _stream_conv2d_4_source_34_source_ram_rdata = (_stream_conv2d_4_source_34_source_sel == 17)? ram_w32_l128_id5_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1333;
  assign stream_conv2d_4_source_34_data = __variable_wdata_1333;
  reg [32-1:0] _stream_conv2d_4_source_34_source_pat_fsm_16;
  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_34_source_pat_all_offset;
  assign _stream_conv2d_4_source_34_source_pat_all_offset = _stream_conv2d_4_source_34_source_offset_buf + _source_stream_conv2d_4_source_34_pat_cur_offset_0 + _source_stream_conv2d_4_source_34_pat_cur_offset_1 + _source_stream_conv2d_4_source_34_pat_cur_offset_2 + _source_stream_conv2d_4_source_34_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_3;
  wire _set_flag_340;
  assign _set_flag_340 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id6_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? _stream_conv2d_4_source_35_source_ram_raddr : 'hx;
  assign ram_w32_l128_id6_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_341 = 1;
  wire [_tmp_341-1:0] _tmp_342;
  assign _tmp_342 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18);
  reg [_tmp_341-1:0] __tmp_342_1;
  assign _stream_conv2d_4_source_35_source_ram_rdata = (_stream_conv2d_4_source_35_source_sel == 18)? ram_w32_l128_id6_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1334;
  assign stream_conv2d_4_source_35_data = __variable_wdata_1334;
  reg [32-1:0] _stream_conv2d_4_source_35_source_pat_fsm_17;
  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_35_source_pat_all_offset;
  assign _stream_conv2d_4_source_35_source_pat_all_offset = _stream_conv2d_4_source_35_source_offset_buf + _source_stream_conv2d_4_source_35_pat_cur_offset_0 + _source_stream_conv2d_4_source_35_pat_cur_offset_1 + _source_stream_conv2d_4_source_35_pat_cur_offset_2 + _source_stream_conv2d_4_source_35_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_3;
  wire _set_flag_343;
  assign _set_flag_343 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id7_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? _stream_conv2d_4_source_36_source_ram_raddr : 'hx;
  assign ram_w32_l128_id7_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_344 = 1;
  wire [_tmp_344-1:0] _tmp_345;
  assign _tmp_345 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19);
  reg [_tmp_344-1:0] __tmp_345_1;
  assign _stream_conv2d_4_source_36_source_ram_rdata = (_stream_conv2d_4_source_36_source_sel == 19)? ram_w32_l128_id7_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1335;
  assign stream_conv2d_4_source_36_data = __variable_wdata_1335;
  reg [32-1:0] _stream_conv2d_4_source_36_source_pat_fsm_18;
  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_36_source_pat_all_offset;
  assign _stream_conv2d_4_source_36_source_pat_all_offset = _stream_conv2d_4_source_36_source_offset_buf + _source_stream_conv2d_4_source_36_pat_cur_offset_0 + _source_stream_conv2d_4_source_36_pat_cur_offset_1 + _source_stream_conv2d_4_source_36_pat_cur_offset_2 + _source_stream_conv2d_4_source_36_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_3;
  wire _set_flag_346;
  assign _set_flag_346 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id8_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? _stream_conv2d_4_source_37_source_ram_raddr : 'hx;
  assign ram_w32_l128_id8_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_347 = 1;
  wire [_tmp_347-1:0] _tmp_348;
  assign _tmp_348 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20);
  reg [_tmp_347-1:0] __tmp_348_1;
  assign _stream_conv2d_4_source_37_source_ram_rdata = (_stream_conv2d_4_source_37_source_sel == 20)? ram_w32_l128_id8_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1336;
  assign stream_conv2d_4_source_37_data = __variable_wdata_1336;
  reg [32-1:0] _stream_conv2d_4_source_37_source_pat_fsm_19;
  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_37_source_pat_all_offset;
  assign _stream_conv2d_4_source_37_source_pat_all_offset = _stream_conv2d_4_source_37_source_offset_buf + _source_stream_conv2d_4_source_37_pat_cur_offset_0 + _source_stream_conv2d_4_source_37_pat_cur_offset_1 + _source_stream_conv2d_4_source_37_pat_cur_offset_2 + _source_stream_conv2d_4_source_37_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_38_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_38_pat_stride_buf_3;
  wire _set_flag_349;
  assign _set_flag_349 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id9_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_38_source_ram_renable && (_stream_conv2d_4_source_38_source_sel == 21))? _stream_conv2d_4_source_38_source_ram_raddr : 'hx;
  assign ram_w32_l128_id9_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_38_source_ram_renable && (_stream_conv2d_4_source_38_source_sel == 21))? 1'd1 : 0;
  localparam _tmp_350 = 1;
  wire [_tmp_350-1:0] _tmp_351;
  assign _tmp_351 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_38_source_ram_renable && (_stream_conv2d_4_source_38_source_sel == 21);
  reg [_tmp_350-1:0] __tmp_351_1;
  assign _stream_conv2d_4_source_38_source_ram_rdata = (_stream_conv2d_4_source_38_source_sel == 21)? ram_w32_l128_id9_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1337;
  assign stream_conv2d_4_source_38_data = __variable_wdata_1337;
  reg [32-1:0] _stream_conv2d_4_source_38_source_pat_fsm_20;
  localparam _stream_conv2d_4_source_38_source_pat_fsm_20_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_38_source_pat_all_offset;
  assign _stream_conv2d_4_source_38_source_pat_all_offset = _stream_conv2d_4_source_38_source_offset_buf + _source_stream_conv2d_4_source_38_pat_cur_offset_0 + _source_stream_conv2d_4_source_38_pat_cur_offset_1 + _source_stream_conv2d_4_source_38_pat_cur_offset_2 + _source_stream_conv2d_4_source_38_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_39_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_39_pat_stride_buf_3;
  wire _set_flag_352;
  assign _set_flag_352 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id10_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_39_source_ram_renable && (_stream_conv2d_4_source_39_source_sel == 22))? _stream_conv2d_4_source_39_source_ram_raddr : 'hx;
  assign ram_w32_l128_id10_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_39_source_ram_renable && (_stream_conv2d_4_source_39_source_sel == 22))? 1'd1 : 0;
  localparam _tmp_353 = 1;
  wire [_tmp_353-1:0] _tmp_354;
  assign _tmp_354 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_39_source_ram_renable && (_stream_conv2d_4_source_39_source_sel == 22);
  reg [_tmp_353-1:0] __tmp_354_1;
  assign _stream_conv2d_4_source_39_source_ram_rdata = (_stream_conv2d_4_source_39_source_sel == 22)? ram_w32_l128_id10_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1338;
  assign stream_conv2d_4_source_39_data = __variable_wdata_1338;
  reg [32-1:0] _stream_conv2d_4_source_39_source_pat_fsm_21;
  localparam _stream_conv2d_4_source_39_source_pat_fsm_21_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_39_source_pat_all_offset;
  assign _stream_conv2d_4_source_39_source_pat_all_offset = _stream_conv2d_4_source_39_source_offset_buf + _source_stream_conv2d_4_source_39_pat_cur_offset_0 + _source_stream_conv2d_4_source_39_pat_cur_offset_1 + _source_stream_conv2d_4_source_39_pat_cur_offset_2 + _source_stream_conv2d_4_source_39_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_40_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_40_pat_stride_buf_3;
  wire _set_flag_355;
  assign _set_flag_355 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id11_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_40_source_ram_renable && (_stream_conv2d_4_source_40_source_sel == 23))? _stream_conv2d_4_source_40_source_ram_raddr : 'hx;
  assign ram_w32_l128_id11_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_40_source_ram_renable && (_stream_conv2d_4_source_40_source_sel == 23))? 1'd1 : 0;
  localparam _tmp_356 = 1;
  wire [_tmp_356-1:0] _tmp_357;
  assign _tmp_357 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_40_source_ram_renable && (_stream_conv2d_4_source_40_source_sel == 23);
  reg [_tmp_356-1:0] __tmp_357_1;
  assign _stream_conv2d_4_source_40_source_ram_rdata = (_stream_conv2d_4_source_40_source_sel == 23)? ram_w32_l128_id11_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1339;
  assign stream_conv2d_4_source_40_data = __variable_wdata_1339;
  reg [32-1:0] _stream_conv2d_4_source_40_source_pat_fsm_22;
  localparam _stream_conv2d_4_source_40_source_pat_fsm_22_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_40_source_pat_all_offset;
  assign _stream_conv2d_4_source_40_source_pat_all_offset = _stream_conv2d_4_source_40_source_offset_buf + _source_stream_conv2d_4_source_40_pat_cur_offset_0 + _source_stream_conv2d_4_source_40_pat_cur_offset_1 + _source_stream_conv2d_4_source_40_pat_cur_offset_2 + _source_stream_conv2d_4_source_40_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_41_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_41_pat_stride_buf_3;
  wire _set_flag_358;
  assign _set_flag_358 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id12_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_41_source_ram_renable && (_stream_conv2d_4_source_41_source_sel == 24))? _stream_conv2d_4_source_41_source_ram_raddr : 'hx;
  assign ram_w32_l128_id12_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_41_source_ram_renable && (_stream_conv2d_4_source_41_source_sel == 24))? 1'd1 : 0;
  localparam _tmp_359 = 1;
  wire [_tmp_359-1:0] _tmp_360;
  assign _tmp_360 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_41_source_ram_renable && (_stream_conv2d_4_source_41_source_sel == 24);
  reg [_tmp_359-1:0] __tmp_360_1;
  assign _stream_conv2d_4_source_41_source_ram_rdata = (_stream_conv2d_4_source_41_source_sel == 24)? ram_w32_l128_id12_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1340;
  assign stream_conv2d_4_source_41_data = __variable_wdata_1340;
  reg [32-1:0] _stream_conv2d_4_source_41_source_pat_fsm_23;
  localparam _stream_conv2d_4_source_41_source_pat_fsm_23_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_41_source_pat_all_offset;
  assign _stream_conv2d_4_source_41_source_pat_all_offset = _stream_conv2d_4_source_41_source_offset_buf + _source_stream_conv2d_4_source_41_pat_cur_offset_0 + _source_stream_conv2d_4_source_41_pat_cur_offset_1 + _source_stream_conv2d_4_source_41_pat_cur_offset_2 + _source_stream_conv2d_4_source_41_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_42_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_42_pat_stride_buf_3;
  wire _set_flag_361;
  assign _set_flag_361 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id13_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_42_source_ram_renable && (_stream_conv2d_4_source_42_source_sel == 25))? _stream_conv2d_4_source_42_source_ram_raddr : 'hx;
  assign ram_w32_l128_id13_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_42_source_ram_renable && (_stream_conv2d_4_source_42_source_sel == 25))? 1'd1 : 0;
  localparam _tmp_362 = 1;
  wire [_tmp_362-1:0] _tmp_363;
  assign _tmp_363 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_42_source_ram_renable && (_stream_conv2d_4_source_42_source_sel == 25);
  reg [_tmp_362-1:0] __tmp_363_1;
  assign _stream_conv2d_4_source_42_source_ram_rdata = (_stream_conv2d_4_source_42_source_sel == 25)? ram_w32_l128_id13_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1341;
  assign stream_conv2d_4_source_42_data = __variable_wdata_1341;
  reg [32-1:0] _stream_conv2d_4_source_42_source_pat_fsm_24;
  localparam _stream_conv2d_4_source_42_source_pat_fsm_24_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_42_source_pat_all_offset;
  assign _stream_conv2d_4_source_42_source_pat_all_offset = _stream_conv2d_4_source_42_source_offset_buf + _source_stream_conv2d_4_source_42_pat_cur_offset_0 + _source_stream_conv2d_4_source_42_pat_cur_offset_1 + _source_stream_conv2d_4_source_42_pat_cur_offset_2 + _source_stream_conv2d_4_source_42_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_43_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_43_pat_stride_buf_3;
  wire _set_flag_364;
  assign _set_flag_364 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id14_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_43_source_ram_renable && (_stream_conv2d_4_source_43_source_sel == 26))? _stream_conv2d_4_source_43_source_ram_raddr : 'hx;
  assign ram_w32_l128_id14_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_43_source_ram_renable && (_stream_conv2d_4_source_43_source_sel == 26))? 1'd1 : 0;
  localparam _tmp_365 = 1;
  wire [_tmp_365-1:0] _tmp_366;
  assign _tmp_366 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_43_source_ram_renable && (_stream_conv2d_4_source_43_source_sel == 26);
  reg [_tmp_365-1:0] __tmp_366_1;
  assign _stream_conv2d_4_source_43_source_ram_rdata = (_stream_conv2d_4_source_43_source_sel == 26)? ram_w32_l128_id14_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1342;
  assign stream_conv2d_4_source_43_data = __variable_wdata_1342;
  reg [32-1:0] _stream_conv2d_4_source_43_source_pat_fsm_25;
  localparam _stream_conv2d_4_source_43_source_pat_fsm_25_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_43_source_pat_all_offset;
  assign _stream_conv2d_4_source_43_source_pat_all_offset = _stream_conv2d_4_source_43_source_offset_buf + _source_stream_conv2d_4_source_43_pat_cur_offset_0 + _source_stream_conv2d_4_source_43_pat_cur_offset_1 + _source_stream_conv2d_4_source_43_pat_cur_offset_2 + _source_stream_conv2d_4_source_43_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_44_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_44_pat_stride_buf_3;
  wire _set_flag_367;
  assign _set_flag_367 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id15_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_44_source_ram_renable && (_stream_conv2d_4_source_44_source_sel == 27))? _stream_conv2d_4_source_44_source_ram_raddr : 'hx;
  assign ram_w32_l128_id15_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_44_source_ram_renable && (_stream_conv2d_4_source_44_source_sel == 27))? 1'd1 : 0;
  localparam _tmp_368 = 1;
  wire [_tmp_368-1:0] _tmp_369;
  assign _tmp_369 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_44_source_ram_renable && (_stream_conv2d_4_source_44_source_sel == 27);
  reg [_tmp_368-1:0] __tmp_369_1;
  assign _stream_conv2d_4_source_44_source_ram_rdata = (_stream_conv2d_4_source_44_source_sel == 27)? ram_w32_l128_id15_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1343;
  assign stream_conv2d_4_source_44_data = __variable_wdata_1343;
  reg [32-1:0] _stream_conv2d_4_source_44_source_pat_fsm_26;
  localparam _stream_conv2d_4_source_44_source_pat_fsm_26_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_44_source_pat_all_offset;
  assign _stream_conv2d_4_source_44_source_pat_all_offset = _stream_conv2d_4_source_44_source_offset_buf + _source_stream_conv2d_4_source_44_pat_cur_offset_0 + _source_stream_conv2d_4_source_44_pat_cur_offset_1 + _source_stream_conv2d_4_source_44_pat_cur_offset_2 + _source_stream_conv2d_4_source_44_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_45_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_45_pat_stride_buf_3;
  wire _set_flag_370;
  assign _set_flag_370 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id16_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_45_source_ram_renable && (_stream_conv2d_4_source_45_source_sel == 28))? _stream_conv2d_4_source_45_source_ram_raddr : 'hx;
  assign ram_w32_l128_id16_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_45_source_ram_renable && (_stream_conv2d_4_source_45_source_sel == 28))? 1'd1 : 0;
  localparam _tmp_371 = 1;
  wire [_tmp_371-1:0] _tmp_372;
  assign _tmp_372 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_45_source_ram_renable && (_stream_conv2d_4_source_45_source_sel == 28);
  reg [_tmp_371-1:0] __tmp_372_1;
  assign _stream_conv2d_4_source_45_source_ram_rdata = (_stream_conv2d_4_source_45_source_sel == 28)? ram_w32_l128_id16_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1344;
  assign stream_conv2d_4_source_45_data = __variable_wdata_1344;
  reg [32-1:0] _stream_conv2d_4_source_45_source_pat_fsm_27;
  localparam _stream_conv2d_4_source_45_source_pat_fsm_27_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_45_source_pat_all_offset;
  assign _stream_conv2d_4_source_45_source_pat_all_offset = _stream_conv2d_4_source_45_source_offset_buf + _source_stream_conv2d_4_source_45_pat_cur_offset_0 + _source_stream_conv2d_4_source_45_pat_cur_offset_1 + _source_stream_conv2d_4_source_45_pat_cur_offset_2 + _source_stream_conv2d_4_source_45_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_46_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_46_pat_stride_buf_3;
  wire _set_flag_373;
  assign _set_flag_373 = conv2d_4_comp_fsm == 3;
  assign ram_w32_l128_id17_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_46_source_ram_renable && (_stream_conv2d_4_source_46_source_sel == 29))? _stream_conv2d_4_source_46_source_ram_raddr : 'hx;
  assign ram_w32_l128_id17_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_46_source_ram_renable && (_stream_conv2d_4_source_46_source_sel == 29))? 1'd1 : 0;
  localparam _tmp_374 = 1;
  wire [_tmp_374-1:0] _tmp_375;
  assign _tmp_375 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_46_source_ram_renable && (_stream_conv2d_4_source_46_source_sel == 29);
  reg [_tmp_374-1:0] __tmp_375_1;
  assign _stream_conv2d_4_source_46_source_ram_rdata = (_stream_conv2d_4_source_46_source_sel == 29)? ram_w32_l128_id17_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_1345;
  assign stream_conv2d_4_source_46_data = __variable_wdata_1345;
  reg [32-1:0] _stream_conv2d_4_source_46_source_pat_fsm_28;
  localparam _stream_conv2d_4_source_46_source_pat_fsm_28_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_46_source_pat_all_offset;
  assign _stream_conv2d_4_source_46_source_pat_all_offset = _stream_conv2d_4_source_46_source_offset_buf + _source_stream_conv2d_4_source_46_pat_cur_offset_0 + _source_stream_conv2d_4_source_46_pat_cur_offset_1 + _source_stream_conv2d_4_source_46_pat_cur_offset_2 + _source_stream_conv2d_4_source_46_pat_cur_offset_3;
  wire _set_flag_376;
  assign _set_flag_376 = conv2d_4_comp_fsm == 3;
  reg _tmp_377;
  reg _tmp_378;
  reg _tmp_379;
  reg _tmp_380;
  reg _tmp_381;
  reg _tmp_382;
  reg _tmp_383;
  reg _tmp_384;
  reg _tmp_385;
  reg _tmp_386;
  reg _tmp_387;
  reg _tmp_388;
  reg _tmp_389;
  reg _tmp_390;
  reg _tmp_391;
  reg _tmp_392;
  reg _tmp_393;
  reg _tmp_394;
  reg _tmp_395;
  reg _tmp_396;
  reg _tmp_397;
  reg _tmp_398;
  reg _tmp_399;
  reg _tmp_400;
  reg _tmp_401;
  reg _tmp_402;
  reg _tmp_403;
  reg _tmp_404;
  reg _tmp_405;
  reg _tmp_406;
  reg _tmp_407;
  reg _tmp_408;
  reg _tmp_409;
  reg _tmp_410;
  reg _tmp_411;
  reg _tmp_412;
  localparam _tmp_413 = 33;
  wire [_tmp_413-1:0] _tmp_414;
  assign _tmp_414 = conv2d_4_stream_out_local + conv2d_4_out_page_comp_offset_buf;
  reg [_tmp_413-1:0] _tmp_415;
  reg [_tmp_413-1:0] _tmp_416;
  reg [_tmp_413-1:0] _tmp_417;
  reg [_tmp_413-1:0] _tmp_418;
  reg [_tmp_413-1:0] _tmp_419;
  reg [_tmp_413-1:0] _tmp_420;
  reg [_tmp_413-1:0] _tmp_421;
  reg [_tmp_413-1:0] _tmp_422;
  reg [_tmp_413-1:0] _tmp_423;
  reg [_tmp_413-1:0] _tmp_424;
  reg [_tmp_413-1:0] _tmp_425;
  reg [_tmp_413-1:0] _tmp_426;
  reg [_tmp_413-1:0] _tmp_427;
  reg [_tmp_413-1:0] _tmp_428;
  reg [_tmp_413-1:0] _tmp_429;
  reg [_tmp_413-1:0] _tmp_430;
  reg [_tmp_413-1:0] _tmp_431;
  reg [_tmp_413-1:0] _tmp_432;
  reg [_tmp_413-1:0] _tmp_433;
  reg [_tmp_413-1:0] _tmp_434;
  reg [_tmp_413-1:0] _tmp_435;
  reg [_tmp_413-1:0] _tmp_436;
  reg [_tmp_413-1:0] _tmp_437;
  reg [_tmp_413-1:0] _tmp_438;
  reg [_tmp_413-1:0] _tmp_439;
  reg [_tmp_413-1:0] _tmp_440;
  reg [_tmp_413-1:0] _tmp_441;
  reg [_tmp_413-1:0] _tmp_442;
  reg [_tmp_413-1:0] _tmp_443;
  reg [_tmp_413-1:0] _tmp_444;
  reg [_tmp_413-1:0] _tmp_445;
  reg [_tmp_413-1:0] _tmp_446;
  reg [_tmp_413-1:0] _tmp_447;
  reg [_tmp_413-1:0] _tmp_448;
  reg [_tmp_413-1:0] _tmp_449;
  reg [_tmp_413-1:0] _tmp_450;
  reg [32-1:0] _tmp_451;
  reg [32-1:0] _tmp_452;
  reg [32-1:0] _tmp_453;
  reg [32-1:0] _tmp_454;
  reg [32-1:0] _tmp_455;
  reg [32-1:0] _tmp_456;
  reg [32-1:0] _tmp_457;
  reg [32-1:0] _tmp_458;
  reg [32-1:0] _tmp_459;
  reg [32-1:0] _tmp_460;
  reg [32-1:0] _tmp_461;
  reg [32-1:0] _tmp_462;
  reg [32-1:0] _tmp_463;
  reg [32-1:0] _tmp_464;
  reg [32-1:0] _tmp_465;
  reg [32-1:0] _tmp_466;
  reg [32-1:0] _tmp_467;
  reg [32-1:0] _tmp_468;
  reg [32-1:0] _tmp_469;
  reg [32-1:0] _tmp_470;
  reg [32-1:0] _tmp_471;
  reg [32-1:0] _tmp_472;
  reg [32-1:0] _tmp_473;
  reg [32-1:0] _tmp_474;
  reg [32-1:0] _tmp_475;
  reg [32-1:0] _tmp_476;
  reg [32-1:0] _tmp_477;
  reg [32-1:0] _tmp_478;
  reg [32-1:0] _tmp_479;
  reg [32-1:0] _tmp_480;
  reg [32-1:0] _tmp_481;
  reg [32-1:0] _tmp_482;
  reg [32-1:0] _tmp_483;
  reg [32-1:0] _tmp_484;
  reg [32-1:0] _tmp_485;
  reg [32-1:0] _tmp_486;
  assign ram_w32_l128_id20_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_89_sink_wenable && (_stream_conv2d_4_sink_89_sink_sel == 30))? _stream_conv2d_4_sink_89_sink_waddr : 'hx;
  assign ram_w32_l128_id20_0_wdata = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_89_sink_wenable && (_stream_conv2d_4_sink_89_sink_sel == 30))? _stream_conv2d_4_sink_89_sink_wdata : 'hx;
  assign ram_w32_l128_id20_0_wenable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_89_sink_wenable && (_stream_conv2d_4_sink_89_sink_sel == 30))? 1'd1 : 0;
  assign ram_w32_l128_id20_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_89_sink_wenable && (_stream_conv2d_4_sink_89_sink_sel == 30))? 1'd1 : 0;
  reg [32-1:0] _stream_conv2d_4_sink_89_sink_fsm_29;
  localparam _stream_conv2d_4_sink_89_sink_fsm_29_init = 0;
  wire _set_flag_487;
  assign _set_flag_487 = conv2d_4_comp_fsm == 4;
  assign _stream_conv2d_4_run_flag = (_set_flag_487)? 1 : 0;
  reg _tmp_488;
  reg _tmp_489;
  reg _tmp_490;
  assign _mul_8_source_stop = _mul_8_stream_oready && 1'd0;
  reg _tmp_491;
  reg _tmp_492;
  reg _tmp_493;
  reg _tmp_494;
  reg _tmp_495;
  reg _tmp_496;
  reg _tmp_497;
  reg _tmp_498;
  reg _tmp_499;
  reg _tmp_500;
  assign _mul_8_sink_start = _tmp_500;
  reg _tmp_501;
  reg _tmp_502;
  reg _tmp_503;
  reg _tmp_504;
  reg _tmp_505;
  reg _tmp_506;
  reg _tmp_507;
  reg _tmp_508;
  reg _tmp_509;
  reg _tmp_510;
  assign _mul_8_sink_stop = _tmp_510;
  reg _tmp_511;
  reg _tmp_512;
  reg _tmp_513;
  reg _tmp_514;
  reg _tmp_515;
  reg _tmp_516;
  reg _tmp_517;
  reg _tmp_518;
  reg _tmp_519;
  reg _tmp_520;
  assign _mul_8_sink_busy = _tmp_520;
  reg _tmp_521;
  assign _mul_8_busy = _mul_8_source_busy || _mul_8_sink_busy || _mul_8_busy_reg;
  reg _tmp_522;
  reg _tmp_523;
  reg _tmp_524;
  assign _mul_9_source_stop = _mul_9_stream_oready && 1'd0;
  reg _tmp_525;
  reg _tmp_526;
  reg _tmp_527;
  reg _tmp_528;
  reg _tmp_529;
  reg _tmp_530;
  reg _tmp_531;
  reg _tmp_532;
  reg _tmp_533;
  reg _tmp_534;
  assign _mul_9_sink_start = _tmp_534;
  reg _tmp_535;
  reg _tmp_536;
  reg _tmp_537;
  reg _tmp_538;
  reg _tmp_539;
  reg _tmp_540;
  reg _tmp_541;
  reg _tmp_542;
  reg _tmp_543;
  reg _tmp_544;
  assign _mul_9_sink_stop = _tmp_544;
  reg _tmp_545;
  reg _tmp_546;
  reg _tmp_547;
  reg _tmp_548;
  reg _tmp_549;
  reg _tmp_550;
  reg _tmp_551;
  reg _tmp_552;
  reg _tmp_553;
  reg _tmp_554;
  assign _mul_9_sink_busy = _tmp_554;
  reg _tmp_555;
  assign _mul_9_busy = _mul_9_source_busy || _mul_9_sink_busy || _mul_9_busy_reg;
  reg _tmp_556;
  reg _tmp_557;
  reg _tmp_558;
  assign _mul_10_source_stop = _mul_10_stream_oready && 1'd0;
  reg _tmp_559;
  reg _tmp_560;
  reg _tmp_561;
  reg _tmp_562;
  reg _tmp_563;
  reg _tmp_564;
  reg _tmp_565;
  reg _tmp_566;
  reg _tmp_567;
  reg _tmp_568;
  assign _mul_10_sink_start = _tmp_568;
  reg _tmp_569;
  reg _tmp_570;
  reg _tmp_571;
  reg _tmp_572;
  reg _tmp_573;
  reg _tmp_574;
  reg _tmp_575;
  reg _tmp_576;
  reg _tmp_577;
  reg _tmp_578;
  assign _mul_10_sink_stop = _tmp_578;
  reg _tmp_579;
  reg _tmp_580;
  reg _tmp_581;
  reg _tmp_582;
  reg _tmp_583;
  reg _tmp_584;
  reg _tmp_585;
  reg _tmp_586;
  reg _tmp_587;
  reg _tmp_588;
  assign _mul_10_sink_busy = _tmp_588;
  reg _tmp_589;
  assign _mul_10_busy = _mul_10_source_busy || _mul_10_sink_busy || _mul_10_busy_reg;
  reg _tmp_590;
  reg _tmp_591;
  reg _tmp_592;
  assign _mul_11_source_stop = _mul_11_stream_oready && 1'd0;
  reg _tmp_593;
  reg _tmp_594;
  reg _tmp_595;
  reg _tmp_596;
  reg _tmp_597;
  reg _tmp_598;
  reg _tmp_599;
  reg _tmp_600;
  reg _tmp_601;
  reg _tmp_602;
  assign _mul_11_sink_start = _tmp_602;
  reg _tmp_603;
  reg _tmp_604;
  reg _tmp_605;
  reg _tmp_606;
  reg _tmp_607;
  reg _tmp_608;
  reg _tmp_609;
  reg _tmp_610;
  reg _tmp_611;
  reg _tmp_612;
  assign _mul_11_sink_stop = _tmp_612;
  reg _tmp_613;
  reg _tmp_614;
  reg _tmp_615;
  reg _tmp_616;
  reg _tmp_617;
  reg _tmp_618;
  reg _tmp_619;
  reg _tmp_620;
  reg _tmp_621;
  reg _tmp_622;
  assign _mul_11_sink_busy = _tmp_622;
  reg _tmp_623;
  assign _mul_11_busy = _mul_11_source_busy || _mul_11_sink_busy || _mul_11_busy_reg;
  reg _tmp_624;
  reg _tmp_625;
  reg _tmp_626;
  assign _mul_12_source_stop = _mul_12_stream_oready && 1'd0;
  reg _tmp_627;
  reg _tmp_628;
  reg _tmp_629;
  reg _tmp_630;
  reg _tmp_631;
  reg _tmp_632;
  reg _tmp_633;
  reg _tmp_634;
  reg _tmp_635;
  reg _tmp_636;
  assign _mul_12_sink_start = _tmp_636;
  reg _tmp_637;
  reg _tmp_638;
  reg _tmp_639;
  reg _tmp_640;
  reg _tmp_641;
  reg _tmp_642;
  reg _tmp_643;
  reg _tmp_644;
  reg _tmp_645;
  reg _tmp_646;
  assign _mul_12_sink_stop = _tmp_646;
  reg _tmp_647;
  reg _tmp_648;
  reg _tmp_649;
  reg _tmp_650;
  reg _tmp_651;
  reg _tmp_652;
  reg _tmp_653;
  reg _tmp_654;
  reg _tmp_655;
  reg _tmp_656;
  assign _mul_12_sink_busy = _tmp_656;
  reg _tmp_657;
  assign _mul_12_busy = _mul_12_source_busy || _mul_12_sink_busy || _mul_12_busy_reg;
  reg _tmp_658;
  reg _tmp_659;
  reg _tmp_660;
  assign _mul_13_source_stop = _mul_13_stream_oready && 1'd0;
  reg _tmp_661;
  reg _tmp_662;
  reg _tmp_663;
  reg _tmp_664;
  reg _tmp_665;
  reg _tmp_666;
  reg _tmp_667;
  reg _tmp_668;
  reg _tmp_669;
  reg _tmp_670;
  assign _mul_13_sink_start = _tmp_670;
  reg _tmp_671;
  reg _tmp_672;
  reg _tmp_673;
  reg _tmp_674;
  reg _tmp_675;
  reg _tmp_676;
  reg _tmp_677;
  reg _tmp_678;
  reg _tmp_679;
  reg _tmp_680;
  assign _mul_13_sink_stop = _tmp_680;
  reg _tmp_681;
  reg _tmp_682;
  reg _tmp_683;
  reg _tmp_684;
  reg _tmp_685;
  reg _tmp_686;
  reg _tmp_687;
  reg _tmp_688;
  reg _tmp_689;
  reg _tmp_690;
  assign _mul_13_sink_busy = _tmp_690;
  reg _tmp_691;
  assign _mul_13_busy = _mul_13_source_busy || _mul_13_sink_busy || _mul_13_busy_reg;
  reg _tmp_692;
  reg _tmp_693;
  reg _tmp_694;
  assign _mul_14_source_stop = _mul_14_stream_oready && 1'd0;
  reg _tmp_695;
  reg _tmp_696;
  reg _tmp_697;
  reg _tmp_698;
  reg _tmp_699;
  reg _tmp_700;
  reg _tmp_701;
  reg _tmp_702;
  reg _tmp_703;
  reg _tmp_704;
  assign _mul_14_sink_start = _tmp_704;
  reg _tmp_705;
  reg _tmp_706;
  reg _tmp_707;
  reg _tmp_708;
  reg _tmp_709;
  reg _tmp_710;
  reg _tmp_711;
  reg _tmp_712;
  reg _tmp_713;
  reg _tmp_714;
  assign _mul_14_sink_stop = _tmp_714;
  reg _tmp_715;
  reg _tmp_716;
  reg _tmp_717;
  reg _tmp_718;
  reg _tmp_719;
  reg _tmp_720;
  reg _tmp_721;
  reg _tmp_722;
  reg _tmp_723;
  reg _tmp_724;
  assign _mul_14_sink_busy = _tmp_724;
  reg _tmp_725;
  assign _mul_14_busy = _mul_14_source_busy || _mul_14_sink_busy || _mul_14_busy_reg;
  reg _tmp_726;
  reg _tmp_727;
  reg _tmp_728;
  assign _mul_15_source_stop = _mul_15_stream_oready && 1'd0;
  reg _tmp_729;
  reg _tmp_730;
  reg _tmp_731;
  reg _tmp_732;
  reg _tmp_733;
  reg _tmp_734;
  reg _tmp_735;
  reg _tmp_736;
  reg _tmp_737;
  reg _tmp_738;
  assign _mul_15_sink_start = _tmp_738;
  reg _tmp_739;
  reg _tmp_740;
  reg _tmp_741;
  reg _tmp_742;
  reg _tmp_743;
  reg _tmp_744;
  reg _tmp_745;
  reg _tmp_746;
  reg _tmp_747;
  reg _tmp_748;
  assign _mul_15_sink_stop = _tmp_748;
  reg _tmp_749;
  reg _tmp_750;
  reg _tmp_751;
  reg _tmp_752;
  reg _tmp_753;
  reg _tmp_754;
  reg _tmp_755;
  reg _tmp_756;
  reg _tmp_757;
  reg _tmp_758;
  assign _mul_15_sink_busy = _tmp_758;
  reg _tmp_759;
  assign _mul_15_busy = _mul_15_source_busy || _mul_15_sink_busy || _mul_15_busy_reg;
  reg _tmp_760;
  reg _tmp_761;
  reg _tmp_762;
  assign _mul_16_source_stop = _mul_16_stream_oready && 1'd0;
  reg _tmp_763;
  reg _tmp_764;
  reg _tmp_765;
  reg _tmp_766;
  reg _tmp_767;
  reg _tmp_768;
  reg _tmp_769;
  reg _tmp_770;
  reg _tmp_771;
  reg _tmp_772;
  assign _mul_16_sink_start = _tmp_772;
  reg _tmp_773;
  reg _tmp_774;
  reg _tmp_775;
  reg _tmp_776;
  reg _tmp_777;
  reg _tmp_778;
  reg _tmp_779;
  reg _tmp_780;
  reg _tmp_781;
  reg _tmp_782;
  assign _mul_16_sink_stop = _tmp_782;
  reg _tmp_783;
  reg _tmp_784;
  reg _tmp_785;
  reg _tmp_786;
  reg _tmp_787;
  reg _tmp_788;
  reg _tmp_789;
  reg _tmp_790;
  reg _tmp_791;
  reg _tmp_792;
  assign _mul_16_sink_busy = _tmp_792;
  reg _tmp_793;
  assign _mul_16_busy = _mul_16_source_busy || _mul_16_sink_busy || _mul_16_busy_reg;
  reg _tmp_794;
  reg _tmp_795;
  reg _tmp_796;
  assign _mul_17_source_stop = _mul_17_stream_oready && 1'd0;
  reg _tmp_797;
  reg _tmp_798;
  reg _tmp_799;
  reg _tmp_800;
  reg _tmp_801;
  reg _tmp_802;
  reg _tmp_803;
  reg _tmp_804;
  reg _tmp_805;
  reg _tmp_806;
  assign _mul_17_sink_start = _tmp_806;
  reg _tmp_807;
  reg _tmp_808;
  reg _tmp_809;
  reg _tmp_810;
  reg _tmp_811;
  reg _tmp_812;
  reg _tmp_813;
  reg _tmp_814;
  reg _tmp_815;
  reg _tmp_816;
  assign _mul_17_sink_stop = _tmp_816;
  reg _tmp_817;
  reg _tmp_818;
  reg _tmp_819;
  reg _tmp_820;
  reg _tmp_821;
  reg _tmp_822;
  reg _tmp_823;
  reg _tmp_824;
  reg _tmp_825;
  reg _tmp_826;
  assign _mul_17_sink_busy = _tmp_826;
  reg _tmp_827;
  assign _mul_17_busy = _mul_17_source_busy || _mul_17_sink_busy || _mul_17_busy_reg;
  reg _tmp_828;
  reg _tmp_829;
  reg _tmp_830;
  assign _mul_18_source_stop = _mul_18_stream_oready && 1'd0;
  reg _tmp_831;
  reg _tmp_832;
  reg _tmp_833;
  reg _tmp_834;
  reg _tmp_835;
  reg _tmp_836;
  reg _tmp_837;
  reg _tmp_838;
  reg _tmp_839;
  reg _tmp_840;
  assign _mul_18_sink_start = _tmp_840;
  reg _tmp_841;
  reg _tmp_842;
  reg _tmp_843;
  reg _tmp_844;
  reg _tmp_845;
  reg _tmp_846;
  reg _tmp_847;
  reg _tmp_848;
  reg _tmp_849;
  reg _tmp_850;
  assign _mul_18_sink_stop = _tmp_850;
  reg _tmp_851;
  reg _tmp_852;
  reg _tmp_853;
  reg _tmp_854;
  reg _tmp_855;
  reg _tmp_856;
  reg _tmp_857;
  reg _tmp_858;
  reg _tmp_859;
  reg _tmp_860;
  assign _mul_18_sink_busy = _tmp_860;
  reg _tmp_861;
  assign _mul_18_busy = _mul_18_source_busy || _mul_18_sink_busy || _mul_18_busy_reg;
  reg _tmp_862;
  reg _tmp_863;
  reg _tmp_864;
  assign _mul_19_source_stop = _mul_19_stream_oready && 1'd0;
  reg _tmp_865;
  reg _tmp_866;
  reg _tmp_867;
  reg _tmp_868;
  reg _tmp_869;
  reg _tmp_870;
  reg _tmp_871;
  reg _tmp_872;
  reg _tmp_873;
  reg _tmp_874;
  assign _mul_19_sink_start = _tmp_874;
  reg _tmp_875;
  reg _tmp_876;
  reg _tmp_877;
  reg _tmp_878;
  reg _tmp_879;
  reg _tmp_880;
  reg _tmp_881;
  reg _tmp_882;
  reg _tmp_883;
  reg _tmp_884;
  assign _mul_19_sink_stop = _tmp_884;
  reg _tmp_885;
  reg _tmp_886;
  reg _tmp_887;
  reg _tmp_888;
  reg _tmp_889;
  reg _tmp_890;
  reg _tmp_891;
  reg _tmp_892;
  reg _tmp_893;
  reg _tmp_894;
  assign _mul_19_sink_busy = _tmp_894;
  reg _tmp_895;
  assign _mul_19_busy = _mul_19_source_busy || _mul_19_sink_busy || _mul_19_busy_reg;
  reg _tmp_896;
  reg _tmp_897;
  reg _tmp_898;
  assign _mul_20_source_stop = _mul_20_stream_oready && 1'd0;
  reg _tmp_899;
  reg _tmp_900;
  reg _tmp_901;
  reg _tmp_902;
  reg _tmp_903;
  reg _tmp_904;
  reg _tmp_905;
  reg _tmp_906;
  reg _tmp_907;
  reg _tmp_908;
  assign _mul_20_sink_start = _tmp_908;
  reg _tmp_909;
  reg _tmp_910;
  reg _tmp_911;
  reg _tmp_912;
  reg _tmp_913;
  reg _tmp_914;
  reg _tmp_915;
  reg _tmp_916;
  reg _tmp_917;
  reg _tmp_918;
  assign _mul_20_sink_stop = _tmp_918;
  reg _tmp_919;
  reg _tmp_920;
  reg _tmp_921;
  reg _tmp_922;
  reg _tmp_923;
  reg _tmp_924;
  reg _tmp_925;
  reg _tmp_926;
  reg _tmp_927;
  reg _tmp_928;
  assign _mul_20_sink_busy = _tmp_928;
  reg _tmp_929;
  assign _mul_20_busy = _mul_20_source_busy || _mul_20_sink_busy || _mul_20_busy_reg;
  reg _tmp_930;
  reg _tmp_931;
  reg _tmp_932;
  assign _mul_21_source_stop = _mul_21_stream_oready && 1'd0;
  reg _tmp_933;
  reg _tmp_934;
  reg _tmp_935;
  reg _tmp_936;
  reg _tmp_937;
  reg _tmp_938;
  reg _tmp_939;
  reg _tmp_940;
  reg _tmp_941;
  reg _tmp_942;
  assign _mul_21_sink_start = _tmp_942;
  reg _tmp_943;
  reg _tmp_944;
  reg _tmp_945;
  reg _tmp_946;
  reg _tmp_947;
  reg _tmp_948;
  reg _tmp_949;
  reg _tmp_950;
  reg _tmp_951;
  reg _tmp_952;
  assign _mul_21_sink_stop = _tmp_952;
  reg _tmp_953;
  reg _tmp_954;
  reg _tmp_955;
  reg _tmp_956;
  reg _tmp_957;
  reg _tmp_958;
  reg _tmp_959;
  reg _tmp_960;
  reg _tmp_961;
  reg _tmp_962;
  assign _mul_21_sink_busy = _tmp_962;
  reg _tmp_963;
  assign _mul_21_busy = _mul_21_source_busy || _mul_21_sink_busy || _mul_21_busy_reg;
  reg _tmp_964;
  reg _tmp_965;
  reg _tmp_966;
  assign _mul_22_source_stop = _mul_22_stream_oready && 1'd0;
  reg _tmp_967;
  reg _tmp_968;
  reg _tmp_969;
  reg _tmp_970;
  reg _tmp_971;
  reg _tmp_972;
  reg _tmp_973;
  reg _tmp_974;
  reg _tmp_975;
  reg _tmp_976;
  assign _mul_22_sink_start = _tmp_976;
  reg _tmp_977;
  reg _tmp_978;
  reg _tmp_979;
  reg _tmp_980;
  reg _tmp_981;
  reg _tmp_982;
  reg _tmp_983;
  reg _tmp_984;
  reg _tmp_985;
  reg _tmp_986;
  assign _mul_22_sink_stop = _tmp_986;
  reg _tmp_987;
  reg _tmp_988;
  reg _tmp_989;
  reg _tmp_990;
  reg _tmp_991;
  reg _tmp_992;
  reg _tmp_993;
  reg _tmp_994;
  reg _tmp_995;
  reg _tmp_996;
  assign _mul_22_sink_busy = _tmp_996;
  reg _tmp_997;
  assign _mul_22_busy = _mul_22_source_busy || _mul_22_sink_busy || _mul_22_busy_reg;
  reg _tmp_998;
  reg _tmp_999;
  reg _tmp_1000;
  assign _mul_23_source_stop = _mul_23_stream_oready && 1'd0;
  reg _tmp_1001;
  reg _tmp_1002;
  reg _tmp_1003;
  reg _tmp_1004;
  reg _tmp_1005;
  reg _tmp_1006;
  reg _tmp_1007;
  reg _tmp_1008;
  reg _tmp_1009;
  reg _tmp_1010;
  assign _mul_23_sink_start = _tmp_1010;
  reg _tmp_1011;
  reg _tmp_1012;
  reg _tmp_1013;
  reg _tmp_1014;
  reg _tmp_1015;
  reg _tmp_1016;
  reg _tmp_1017;
  reg _tmp_1018;
  reg _tmp_1019;
  reg _tmp_1020;
  assign _mul_23_sink_stop = _tmp_1020;
  reg _tmp_1021;
  reg _tmp_1022;
  reg _tmp_1023;
  reg _tmp_1024;
  reg _tmp_1025;
  reg _tmp_1026;
  reg _tmp_1027;
  reg _tmp_1028;
  reg _tmp_1029;
  reg _tmp_1030;
  assign _mul_23_sink_busy = _tmp_1030;
  reg _tmp_1031;
  assign _mul_23_busy = _mul_23_source_busy || _mul_23_sink_busy || _mul_23_busy_reg;
  reg _tmp_1032;
  reg _tmp_1033;
  reg _tmp_1034;
  assign _mul_24_source_stop = _mul_24_stream_oready && 1'd0;
  reg _tmp_1035;
  reg _tmp_1036;
  reg _tmp_1037;
  reg _tmp_1038;
  reg _tmp_1039;
  reg _tmp_1040;
  reg _tmp_1041;
  reg _tmp_1042;
  reg _tmp_1043;
  reg _tmp_1044;
  assign _mul_24_sink_start = _tmp_1044;
  reg _tmp_1045;
  reg _tmp_1046;
  reg _tmp_1047;
  reg _tmp_1048;
  reg _tmp_1049;
  reg _tmp_1050;
  reg _tmp_1051;
  reg _tmp_1052;
  reg _tmp_1053;
  reg _tmp_1054;
  assign _mul_24_sink_stop = _tmp_1054;
  reg _tmp_1055;
  reg _tmp_1056;
  reg _tmp_1057;
  reg _tmp_1058;
  reg _tmp_1059;
  reg _tmp_1060;
  reg _tmp_1061;
  reg _tmp_1062;
  reg _tmp_1063;
  reg _tmp_1064;
  assign _mul_24_sink_busy = _tmp_1064;
  reg _tmp_1065;
  assign _mul_24_busy = _mul_24_source_busy || _mul_24_sink_busy || _mul_24_busy_reg;
  reg _tmp_1066;
  reg _tmp_1067;
  reg _tmp_1068;
  assign _mul_25_source_stop = _mul_25_stream_oready && 1'd0;
  reg _tmp_1069;
  reg _tmp_1070;
  reg _tmp_1071;
  reg _tmp_1072;
  reg _tmp_1073;
  reg _tmp_1074;
  reg _tmp_1075;
  reg _tmp_1076;
  reg _tmp_1077;
  reg _tmp_1078;
  assign _mul_25_sink_start = _tmp_1078;
  reg _tmp_1079;
  reg _tmp_1080;
  reg _tmp_1081;
  reg _tmp_1082;
  reg _tmp_1083;
  reg _tmp_1084;
  reg _tmp_1085;
  reg _tmp_1086;
  reg _tmp_1087;
  reg _tmp_1088;
  assign _mul_25_sink_stop = _tmp_1088;
  reg _tmp_1089;
  reg _tmp_1090;
  reg _tmp_1091;
  reg _tmp_1092;
  reg _tmp_1093;
  reg _tmp_1094;
  reg _tmp_1095;
  reg _tmp_1096;
  reg _tmp_1097;
  reg _tmp_1098;
  assign _mul_25_sink_busy = _tmp_1098;
  reg _tmp_1099;
  assign _mul_25_busy = _mul_25_source_busy || _mul_25_sink_busy || _mul_25_busy_reg;
  reg _tmp_1100;
  reg _tmp_1101;
  reg _tmp_1102;
  assign _add_tree_4_source_stop = _add_tree_4_stream_oready && 1'd0;
  reg _tmp_1103;
  reg _tmp_1104;
  reg _tmp_1105;
  reg _tmp_1106;
  reg _tmp_1107;
  assign _add_tree_4_sink_start = _tmp_1107;
  reg _tmp_1108;
  reg _tmp_1109;
  reg _tmp_1110;
  reg _tmp_1111;
  reg _tmp_1112;
  assign _add_tree_4_sink_stop = _tmp_1112;
  reg _tmp_1113;
  reg _tmp_1114;
  reg _tmp_1115;
  reg _tmp_1116;
  reg _tmp_1117;
  assign _add_tree_4_sink_busy = _tmp_1117;
  reg _tmp_1118;
  assign _add_tree_4_busy = _add_tree_4_source_busy || _add_tree_4_sink_busy || _add_tree_4_busy_reg;
  reg _tmp_1119;
  reg _tmp_1120;
  reg _tmp_1121;
  reg _tmp_1122;
  reg _tmp_1123;
  reg _tmp_1124;
  reg _tmp_1125;
  reg _tmp_1126;
  reg _tmp_1127;
  reg _tmp_1128;
  assign _acc_0_source_stop = _acc_0_stream_oready && 1'd0;
  reg _tmp_1129;
  reg _tmp_1130;
  reg _tmp_1131;
  reg _tmp_1132;
  reg _tmp_1133;
  reg _tmp_1134;
  reg _tmp_1135;
  assign _acc_0_sink_start = _tmp_1135;
  reg _tmp_1136;
  reg _tmp_1137;
  reg _tmp_1138;
  reg _tmp_1139;
  reg _tmp_1140;
  reg _tmp_1141;
  reg _tmp_1142;
  assign _acc_0_sink_stop = _tmp_1142;
  reg _tmp_1143;
  reg _tmp_1144;
  reg _tmp_1145;
  reg _tmp_1146;
  reg _tmp_1147;
  reg _tmp_1148;
  reg _tmp_1149;
  assign _acc_0_sink_busy = _tmp_1149;
  reg _tmp_1150;
  assign _acc_0_busy = _acc_0_source_busy || _acc_0_sink_busy || _acc_0_busy_reg;
  reg _tmp_1151;
  reg _tmp_1152;
  reg _tmp_1153;
  assign _mul_rshift_round_clip_6_source_stop = _mul_rshift_round_clip_6_stream_oready && 1'd0;
  reg _tmp_1154;
  reg _tmp_1155;
  reg _tmp_1156;
  reg _tmp_1157;
  reg _tmp_1158;
  reg _tmp_1159;
  reg _tmp_1160;
  reg _tmp_1161;
  reg _tmp_1162;
  reg _tmp_1163;
  assign _mul_rshift_round_clip_6_sink_start = _tmp_1163;
  reg _tmp_1164;
  reg _tmp_1165;
  reg _tmp_1166;
  reg _tmp_1167;
  reg _tmp_1168;
  reg _tmp_1169;
  reg _tmp_1170;
  reg _tmp_1171;
  reg _tmp_1172;
  reg _tmp_1173;
  assign _mul_rshift_round_clip_6_sink_stop = _tmp_1173;
  reg _tmp_1174;
  reg _tmp_1175;
  reg _tmp_1176;
  reg _tmp_1177;
  reg _tmp_1178;
  reg _tmp_1179;
  reg _tmp_1180;
  reg _tmp_1181;
  reg _tmp_1182;
  reg _tmp_1183;
  assign _mul_rshift_round_clip_6_sink_busy = _tmp_1183;
  reg _tmp_1184;
  assign _mul_rshift_round_clip_6_busy = _mul_rshift_round_clip_6_source_busy || _mul_rshift_round_clip_6_sink_busy || _mul_rshift_round_clip_6_busy_reg;
  reg _tmp_1185;
  reg _tmp_1186;
  reg _tmp_1187;
  assign _mul_26_source_stop = _mul_26_stream_oready && 1'd0;
  reg _tmp_1188;
  reg _tmp_1189;
  reg _tmp_1190;
  reg _tmp_1191;
  reg _tmp_1192;
  reg _tmp_1193;
  reg _tmp_1194;
  reg _tmp_1195;
  reg _tmp_1196;
  reg _tmp_1197;
  assign _mul_26_sink_start = _tmp_1197;
  reg _tmp_1198;
  reg _tmp_1199;
  reg _tmp_1200;
  reg _tmp_1201;
  reg _tmp_1202;
  reg _tmp_1203;
  reg _tmp_1204;
  reg _tmp_1205;
  reg _tmp_1206;
  reg _tmp_1207;
  assign _mul_26_sink_stop = _tmp_1207;
  reg _tmp_1208;
  reg _tmp_1209;
  reg _tmp_1210;
  reg _tmp_1211;
  reg _tmp_1212;
  reg _tmp_1213;
  reg _tmp_1214;
  reg _tmp_1215;
  reg _tmp_1216;
  reg _tmp_1217;
  assign _mul_26_sink_busy = _tmp_1217;
  reg _tmp_1218;
  assign _mul_26_busy = _mul_26_source_busy || _mul_26_sink_busy || _mul_26_busy_reg;
  reg _tmp_1219;
  reg _tmp_1220;
  reg _tmp_1221;
  assign _mul_27_source_stop = _mul_27_stream_oready && 1'd0;
  reg _tmp_1222;
  reg _tmp_1223;
  reg _tmp_1224;
  reg _tmp_1225;
  reg _tmp_1226;
  reg _tmp_1227;
  reg _tmp_1228;
  reg _tmp_1229;
  reg _tmp_1230;
  reg _tmp_1231;
  assign _mul_27_sink_start = _tmp_1231;
  reg _tmp_1232;
  reg _tmp_1233;
  reg _tmp_1234;
  reg _tmp_1235;
  reg _tmp_1236;
  reg _tmp_1237;
  reg _tmp_1238;
  reg _tmp_1239;
  reg _tmp_1240;
  reg _tmp_1241;
  assign _mul_27_sink_stop = _tmp_1241;
  reg _tmp_1242;
  reg _tmp_1243;
  reg _tmp_1244;
  reg _tmp_1245;
  reg _tmp_1246;
  reg _tmp_1247;
  reg _tmp_1248;
  reg _tmp_1249;
  reg _tmp_1250;
  reg _tmp_1251;
  assign _mul_27_sink_busy = _tmp_1251;
  reg _tmp_1252;
  assign _mul_27_busy = _mul_27_source_busy || _mul_27_sink_busy || _mul_27_busy_reg;
  reg _tmp_1253;
  reg _tmp_1254;
  reg _tmp_1255;
  assign _mul_28_source_stop = _mul_28_stream_oready && 1'd0;
  reg _tmp_1256;
  reg _tmp_1257;
  reg _tmp_1258;
  reg _tmp_1259;
  reg _tmp_1260;
  reg _tmp_1261;
  reg _tmp_1262;
  reg _tmp_1263;
  reg _tmp_1264;
  reg _tmp_1265;
  assign _mul_28_sink_start = _tmp_1265;
  reg _tmp_1266;
  reg _tmp_1267;
  reg _tmp_1268;
  reg _tmp_1269;
  reg _tmp_1270;
  reg _tmp_1271;
  reg _tmp_1272;
  reg _tmp_1273;
  reg _tmp_1274;
  reg _tmp_1275;
  assign _mul_28_sink_stop = _tmp_1275;
  reg _tmp_1276;
  reg _tmp_1277;
  reg _tmp_1278;
  reg _tmp_1279;
  reg _tmp_1280;
  reg _tmp_1281;
  reg _tmp_1282;
  reg _tmp_1283;
  reg _tmp_1284;
  reg _tmp_1285;
  assign _mul_28_sink_busy = _tmp_1285;
  reg _tmp_1286;
  assign _mul_28_busy = _mul_28_source_busy || _mul_28_sink_busy || _mul_28_busy_reg;
  reg _tmp_1287;
  reg _tmp_1288;
  reg _tmp_1289;
  assign _mul_29_source_stop = _mul_29_stream_oready && 1'd0;
  reg _tmp_1290;
  reg _tmp_1291;
  reg _tmp_1292;
  reg _tmp_1293;
  reg _tmp_1294;
  reg _tmp_1295;
  reg _tmp_1296;
  reg _tmp_1297;
  reg _tmp_1298;
  reg _tmp_1299;
  assign _mul_29_sink_start = _tmp_1299;
  reg _tmp_1300;
  reg _tmp_1301;
  reg _tmp_1302;
  reg _tmp_1303;
  reg _tmp_1304;
  reg _tmp_1305;
  reg _tmp_1306;
  reg _tmp_1307;
  reg _tmp_1308;
  reg _tmp_1309;
  assign _mul_29_sink_stop = _tmp_1309;
  reg _tmp_1310;
  reg _tmp_1311;
  reg _tmp_1312;
  reg _tmp_1313;
  reg _tmp_1314;
  reg _tmp_1315;
  reg _tmp_1316;
  reg _tmp_1317;
  reg _tmp_1318;
  reg _tmp_1319;
  assign _mul_29_sink_busy = _tmp_1319;
  reg _tmp_1320;
  assign _mul_29_busy = _mul_29_source_busy || _mul_29_sink_busy || _mul_29_busy_reg;
  reg _tmp_1321;
  reg _tmp_1322;
  reg _tmp_1323;
  assign _mul_30_source_stop = _mul_30_stream_oready && 1'd0;
  reg _tmp_1324;
  reg _tmp_1325;
  reg _tmp_1326;
  reg _tmp_1327;
  reg _tmp_1328;
  reg _tmp_1329;
  reg _tmp_1330;
  reg _tmp_1331;
  reg _tmp_1332;
  reg _tmp_1333;
  assign _mul_30_sink_start = _tmp_1333;
  reg _tmp_1334;
  reg _tmp_1335;
  reg _tmp_1336;
  reg _tmp_1337;
  reg _tmp_1338;
  reg _tmp_1339;
  reg _tmp_1340;
  reg _tmp_1341;
  reg _tmp_1342;
  reg _tmp_1343;
  assign _mul_30_sink_stop = _tmp_1343;
  reg _tmp_1344;
  reg _tmp_1345;
  reg _tmp_1346;
  reg _tmp_1347;
  reg _tmp_1348;
  reg _tmp_1349;
  reg _tmp_1350;
  reg _tmp_1351;
  reg _tmp_1352;
  reg _tmp_1353;
  assign _mul_30_sink_busy = _tmp_1353;
  reg _tmp_1354;
  assign _mul_30_busy = _mul_30_source_busy || _mul_30_sink_busy || _mul_30_busy_reg;
  reg _tmp_1355;
  reg _tmp_1356;
  reg _tmp_1357;
  assign _mul_31_source_stop = _mul_31_stream_oready && 1'd0;
  reg _tmp_1358;
  reg _tmp_1359;
  reg _tmp_1360;
  reg _tmp_1361;
  reg _tmp_1362;
  reg _tmp_1363;
  reg _tmp_1364;
  reg _tmp_1365;
  reg _tmp_1366;
  reg _tmp_1367;
  assign _mul_31_sink_start = _tmp_1367;
  reg _tmp_1368;
  reg _tmp_1369;
  reg _tmp_1370;
  reg _tmp_1371;
  reg _tmp_1372;
  reg _tmp_1373;
  reg _tmp_1374;
  reg _tmp_1375;
  reg _tmp_1376;
  reg _tmp_1377;
  assign _mul_31_sink_stop = _tmp_1377;
  reg _tmp_1378;
  reg _tmp_1379;
  reg _tmp_1380;
  reg _tmp_1381;
  reg _tmp_1382;
  reg _tmp_1383;
  reg _tmp_1384;
  reg _tmp_1385;
  reg _tmp_1386;
  reg _tmp_1387;
  assign _mul_31_sink_busy = _tmp_1387;
  reg _tmp_1388;
  assign _mul_31_busy = _mul_31_source_busy || _mul_31_sink_busy || _mul_31_busy_reg;
  reg _tmp_1389;
  reg _tmp_1390;
  reg _tmp_1391;
  assign _mul_32_source_stop = _mul_32_stream_oready && 1'd0;
  reg _tmp_1392;
  reg _tmp_1393;
  reg _tmp_1394;
  reg _tmp_1395;
  reg _tmp_1396;
  reg _tmp_1397;
  reg _tmp_1398;
  reg _tmp_1399;
  reg _tmp_1400;
  reg _tmp_1401;
  assign _mul_32_sink_start = _tmp_1401;
  reg _tmp_1402;
  reg _tmp_1403;
  reg _tmp_1404;
  reg _tmp_1405;
  reg _tmp_1406;
  reg _tmp_1407;
  reg _tmp_1408;
  reg _tmp_1409;
  reg _tmp_1410;
  reg _tmp_1411;
  assign _mul_32_sink_stop = _tmp_1411;
  reg _tmp_1412;
  reg _tmp_1413;
  reg _tmp_1414;
  reg _tmp_1415;
  reg _tmp_1416;
  reg _tmp_1417;
  reg _tmp_1418;
  reg _tmp_1419;
  reg _tmp_1420;
  reg _tmp_1421;
  assign _mul_32_sink_busy = _tmp_1421;
  reg _tmp_1422;
  assign _mul_32_busy = _mul_32_source_busy || _mul_32_sink_busy || _mul_32_busy_reg;
  reg _tmp_1423;
  reg _tmp_1424;
  reg _tmp_1425;
  assign _mul_33_source_stop = _mul_33_stream_oready && 1'd0;
  reg _tmp_1426;
  reg _tmp_1427;
  reg _tmp_1428;
  reg _tmp_1429;
  reg _tmp_1430;
  reg _tmp_1431;
  reg _tmp_1432;
  reg _tmp_1433;
  reg _tmp_1434;
  reg _tmp_1435;
  assign _mul_33_sink_start = _tmp_1435;
  reg _tmp_1436;
  reg _tmp_1437;
  reg _tmp_1438;
  reg _tmp_1439;
  reg _tmp_1440;
  reg _tmp_1441;
  reg _tmp_1442;
  reg _tmp_1443;
  reg _tmp_1444;
  reg _tmp_1445;
  assign _mul_33_sink_stop = _tmp_1445;
  reg _tmp_1446;
  reg _tmp_1447;
  reg _tmp_1448;
  reg _tmp_1449;
  reg _tmp_1450;
  reg _tmp_1451;
  reg _tmp_1452;
  reg _tmp_1453;
  reg _tmp_1454;
  reg _tmp_1455;
  assign _mul_33_sink_busy = _tmp_1455;
  reg _tmp_1456;
  assign _mul_33_busy = _mul_33_source_busy || _mul_33_sink_busy || _mul_33_busy_reg;
  reg _tmp_1457;
  reg _tmp_1458;
  reg _tmp_1459;
  assign _mul_34_source_stop = _mul_34_stream_oready && 1'd0;
  reg _tmp_1460;
  reg _tmp_1461;
  reg _tmp_1462;
  reg _tmp_1463;
  reg _tmp_1464;
  reg _tmp_1465;
  reg _tmp_1466;
  reg _tmp_1467;
  reg _tmp_1468;
  reg _tmp_1469;
  assign _mul_34_sink_start = _tmp_1469;
  reg _tmp_1470;
  reg _tmp_1471;
  reg _tmp_1472;
  reg _tmp_1473;
  reg _tmp_1474;
  reg _tmp_1475;
  reg _tmp_1476;
  reg _tmp_1477;
  reg _tmp_1478;
  reg _tmp_1479;
  assign _mul_34_sink_stop = _tmp_1479;
  reg _tmp_1480;
  reg _tmp_1481;
  reg _tmp_1482;
  reg _tmp_1483;
  reg _tmp_1484;
  reg _tmp_1485;
  reg _tmp_1486;
  reg _tmp_1487;
  reg _tmp_1488;
  reg _tmp_1489;
  assign _mul_34_sink_busy = _tmp_1489;
  reg _tmp_1490;
  assign _mul_34_busy = _mul_34_source_busy || _mul_34_sink_busy || _mul_34_busy_reg;
  reg _tmp_1491;
  reg _tmp_1492;
  reg _tmp_1493;
  assign _mul_35_source_stop = _mul_35_stream_oready && 1'd0;
  reg _tmp_1494;
  reg _tmp_1495;
  reg _tmp_1496;
  reg _tmp_1497;
  reg _tmp_1498;
  reg _tmp_1499;
  reg _tmp_1500;
  reg _tmp_1501;
  reg _tmp_1502;
  reg _tmp_1503;
  assign _mul_35_sink_start = _tmp_1503;
  reg _tmp_1504;
  reg _tmp_1505;
  reg _tmp_1506;
  reg _tmp_1507;
  reg _tmp_1508;
  reg _tmp_1509;
  reg _tmp_1510;
  reg _tmp_1511;
  reg _tmp_1512;
  reg _tmp_1513;
  assign _mul_35_sink_stop = _tmp_1513;
  reg _tmp_1514;
  reg _tmp_1515;
  reg _tmp_1516;
  reg _tmp_1517;
  reg _tmp_1518;
  reg _tmp_1519;
  reg _tmp_1520;
  reg _tmp_1521;
  reg _tmp_1522;
  reg _tmp_1523;
  assign _mul_35_sink_busy = _tmp_1523;
  reg _tmp_1524;
  assign _mul_35_busy = _mul_35_source_busy || _mul_35_sink_busy || _mul_35_busy_reg;
  reg _tmp_1525;
  reg _tmp_1526;
  reg _tmp_1527;
  assign _mul_36_source_stop = _mul_36_stream_oready && 1'd0;
  reg _tmp_1528;
  reg _tmp_1529;
  reg _tmp_1530;
  reg _tmp_1531;
  reg _tmp_1532;
  reg _tmp_1533;
  reg _tmp_1534;
  reg _tmp_1535;
  reg _tmp_1536;
  reg _tmp_1537;
  assign _mul_36_sink_start = _tmp_1537;
  reg _tmp_1538;
  reg _tmp_1539;
  reg _tmp_1540;
  reg _tmp_1541;
  reg _tmp_1542;
  reg _tmp_1543;
  reg _tmp_1544;
  reg _tmp_1545;
  reg _tmp_1546;
  reg _tmp_1547;
  assign _mul_36_sink_stop = _tmp_1547;
  reg _tmp_1548;
  reg _tmp_1549;
  reg _tmp_1550;
  reg _tmp_1551;
  reg _tmp_1552;
  reg _tmp_1553;
  reg _tmp_1554;
  reg _tmp_1555;
  reg _tmp_1556;
  reg _tmp_1557;
  assign _mul_36_sink_busy = _tmp_1557;
  reg _tmp_1558;
  assign _mul_36_busy = _mul_36_source_busy || _mul_36_sink_busy || _mul_36_busy_reg;
  reg _tmp_1559;
  reg _tmp_1560;
  reg _tmp_1561;
  assign _mul_37_source_stop = _mul_37_stream_oready && 1'd0;
  reg _tmp_1562;
  reg _tmp_1563;
  reg _tmp_1564;
  reg _tmp_1565;
  reg _tmp_1566;
  reg _tmp_1567;
  reg _tmp_1568;
  reg _tmp_1569;
  reg _tmp_1570;
  reg _tmp_1571;
  assign _mul_37_sink_start = _tmp_1571;
  reg _tmp_1572;
  reg _tmp_1573;
  reg _tmp_1574;
  reg _tmp_1575;
  reg _tmp_1576;
  reg _tmp_1577;
  reg _tmp_1578;
  reg _tmp_1579;
  reg _tmp_1580;
  reg _tmp_1581;
  assign _mul_37_sink_stop = _tmp_1581;
  reg _tmp_1582;
  reg _tmp_1583;
  reg _tmp_1584;
  reg _tmp_1585;
  reg _tmp_1586;
  reg _tmp_1587;
  reg _tmp_1588;
  reg _tmp_1589;
  reg _tmp_1590;
  reg _tmp_1591;
  assign _mul_37_sink_busy = _tmp_1591;
  reg _tmp_1592;
  assign _mul_37_busy = _mul_37_source_busy || _mul_37_sink_busy || _mul_37_busy_reg;
  reg _tmp_1593;
  reg _tmp_1594;
  reg _tmp_1595;
  assign _mul_38_source_stop = _mul_38_stream_oready && 1'd0;
  reg _tmp_1596;
  reg _tmp_1597;
  reg _tmp_1598;
  reg _tmp_1599;
  reg _tmp_1600;
  reg _tmp_1601;
  reg _tmp_1602;
  reg _tmp_1603;
  reg _tmp_1604;
  reg _tmp_1605;
  assign _mul_38_sink_start = _tmp_1605;
  reg _tmp_1606;
  reg _tmp_1607;
  reg _tmp_1608;
  reg _tmp_1609;
  reg _tmp_1610;
  reg _tmp_1611;
  reg _tmp_1612;
  reg _tmp_1613;
  reg _tmp_1614;
  reg _tmp_1615;
  assign _mul_38_sink_stop = _tmp_1615;
  reg _tmp_1616;
  reg _tmp_1617;
  reg _tmp_1618;
  reg _tmp_1619;
  reg _tmp_1620;
  reg _tmp_1621;
  reg _tmp_1622;
  reg _tmp_1623;
  reg _tmp_1624;
  reg _tmp_1625;
  assign _mul_38_sink_busy = _tmp_1625;
  reg _tmp_1626;
  assign _mul_38_busy = _mul_38_source_busy || _mul_38_sink_busy || _mul_38_busy_reg;
  reg _tmp_1627;
  reg _tmp_1628;
  reg _tmp_1629;
  assign _mul_39_source_stop = _mul_39_stream_oready && 1'd0;
  reg _tmp_1630;
  reg _tmp_1631;
  reg _tmp_1632;
  reg _tmp_1633;
  reg _tmp_1634;
  reg _tmp_1635;
  reg _tmp_1636;
  reg _tmp_1637;
  reg _tmp_1638;
  reg _tmp_1639;
  assign _mul_39_sink_start = _tmp_1639;
  reg _tmp_1640;
  reg _tmp_1641;
  reg _tmp_1642;
  reg _tmp_1643;
  reg _tmp_1644;
  reg _tmp_1645;
  reg _tmp_1646;
  reg _tmp_1647;
  reg _tmp_1648;
  reg _tmp_1649;
  assign _mul_39_sink_stop = _tmp_1649;
  reg _tmp_1650;
  reg _tmp_1651;
  reg _tmp_1652;
  reg _tmp_1653;
  reg _tmp_1654;
  reg _tmp_1655;
  reg _tmp_1656;
  reg _tmp_1657;
  reg _tmp_1658;
  reg _tmp_1659;
  assign _mul_39_sink_busy = _tmp_1659;
  reg _tmp_1660;
  assign _mul_39_busy = _mul_39_source_busy || _mul_39_sink_busy || _mul_39_busy_reg;
  reg _tmp_1661;
  reg _tmp_1662;
  reg _tmp_1663;
  assign _mul_40_source_stop = _mul_40_stream_oready && 1'd0;
  reg _tmp_1664;
  reg _tmp_1665;
  reg _tmp_1666;
  reg _tmp_1667;
  reg _tmp_1668;
  reg _tmp_1669;
  reg _tmp_1670;
  reg _tmp_1671;
  reg _tmp_1672;
  reg _tmp_1673;
  assign _mul_40_sink_start = _tmp_1673;
  reg _tmp_1674;
  reg _tmp_1675;
  reg _tmp_1676;
  reg _tmp_1677;
  reg _tmp_1678;
  reg _tmp_1679;
  reg _tmp_1680;
  reg _tmp_1681;
  reg _tmp_1682;
  reg _tmp_1683;
  assign _mul_40_sink_stop = _tmp_1683;
  reg _tmp_1684;
  reg _tmp_1685;
  reg _tmp_1686;
  reg _tmp_1687;
  reg _tmp_1688;
  reg _tmp_1689;
  reg _tmp_1690;
  reg _tmp_1691;
  reg _tmp_1692;
  reg _tmp_1693;
  assign _mul_40_sink_busy = _tmp_1693;
  reg _tmp_1694;
  assign _mul_40_busy = _mul_40_source_busy || _mul_40_sink_busy || _mul_40_busy_reg;
  reg _tmp_1695;
  reg _tmp_1696;
  reg _tmp_1697;
  assign _mul_41_source_stop = _mul_41_stream_oready && 1'd0;
  reg _tmp_1698;
  reg _tmp_1699;
  reg _tmp_1700;
  reg _tmp_1701;
  reg _tmp_1702;
  reg _tmp_1703;
  reg _tmp_1704;
  reg _tmp_1705;
  reg _tmp_1706;
  reg _tmp_1707;
  assign _mul_41_sink_start = _tmp_1707;
  reg _tmp_1708;
  reg _tmp_1709;
  reg _tmp_1710;
  reg _tmp_1711;
  reg _tmp_1712;
  reg _tmp_1713;
  reg _tmp_1714;
  reg _tmp_1715;
  reg _tmp_1716;
  reg _tmp_1717;
  assign _mul_41_sink_stop = _tmp_1717;
  reg _tmp_1718;
  reg _tmp_1719;
  reg _tmp_1720;
  reg _tmp_1721;
  reg _tmp_1722;
  reg _tmp_1723;
  reg _tmp_1724;
  reg _tmp_1725;
  reg _tmp_1726;
  reg _tmp_1727;
  assign _mul_41_sink_busy = _tmp_1727;
  reg _tmp_1728;
  assign _mul_41_busy = _mul_41_source_busy || _mul_41_sink_busy || _mul_41_busy_reg;
  reg _tmp_1729;
  reg _tmp_1730;
  reg _tmp_1731;
  assign _mul_42_source_stop = _mul_42_stream_oready && 1'd0;
  reg _tmp_1732;
  reg _tmp_1733;
  reg _tmp_1734;
  reg _tmp_1735;
  reg _tmp_1736;
  reg _tmp_1737;
  reg _tmp_1738;
  reg _tmp_1739;
  reg _tmp_1740;
  reg _tmp_1741;
  assign _mul_42_sink_start = _tmp_1741;
  reg _tmp_1742;
  reg _tmp_1743;
  reg _tmp_1744;
  reg _tmp_1745;
  reg _tmp_1746;
  reg _tmp_1747;
  reg _tmp_1748;
  reg _tmp_1749;
  reg _tmp_1750;
  reg _tmp_1751;
  assign _mul_42_sink_stop = _tmp_1751;
  reg _tmp_1752;
  reg _tmp_1753;
  reg _tmp_1754;
  reg _tmp_1755;
  reg _tmp_1756;
  reg _tmp_1757;
  reg _tmp_1758;
  reg _tmp_1759;
  reg _tmp_1760;
  reg _tmp_1761;
  assign _mul_42_sink_busy = _tmp_1761;
  reg _tmp_1762;
  assign _mul_42_busy = _mul_42_source_busy || _mul_42_sink_busy || _mul_42_busy_reg;
  reg _tmp_1763;
  reg _tmp_1764;
  reg _tmp_1765;
  assign _mul_43_source_stop = _mul_43_stream_oready && 1'd0;
  reg _tmp_1766;
  reg _tmp_1767;
  reg _tmp_1768;
  reg _tmp_1769;
  reg _tmp_1770;
  reg _tmp_1771;
  reg _tmp_1772;
  reg _tmp_1773;
  reg _tmp_1774;
  reg _tmp_1775;
  assign _mul_43_sink_start = _tmp_1775;
  reg _tmp_1776;
  reg _tmp_1777;
  reg _tmp_1778;
  reg _tmp_1779;
  reg _tmp_1780;
  reg _tmp_1781;
  reg _tmp_1782;
  reg _tmp_1783;
  reg _tmp_1784;
  reg _tmp_1785;
  assign _mul_43_sink_stop = _tmp_1785;
  reg _tmp_1786;
  reg _tmp_1787;
  reg _tmp_1788;
  reg _tmp_1789;
  reg _tmp_1790;
  reg _tmp_1791;
  reg _tmp_1792;
  reg _tmp_1793;
  reg _tmp_1794;
  reg _tmp_1795;
  assign _mul_43_sink_busy = _tmp_1795;
  reg _tmp_1796;
  assign _mul_43_busy = _mul_43_source_busy || _mul_43_sink_busy || _mul_43_busy_reg;
  reg _tmp_1797;
  reg _tmp_1798;
  reg _tmp_1799;
  assign _add_tree_5_source_stop = _add_tree_5_stream_oready && 1'd0;
  reg _tmp_1800;
  reg _tmp_1801;
  reg _tmp_1802;
  reg _tmp_1803;
  reg _tmp_1804;
  assign _add_tree_5_sink_start = _tmp_1804;
  reg _tmp_1805;
  reg _tmp_1806;
  reg _tmp_1807;
  reg _tmp_1808;
  reg _tmp_1809;
  assign _add_tree_5_sink_stop = _tmp_1809;
  reg _tmp_1810;
  reg _tmp_1811;
  reg _tmp_1812;
  reg _tmp_1813;
  reg _tmp_1814;
  assign _add_tree_5_sink_busy = _tmp_1814;
  reg _tmp_1815;
  assign _add_tree_5_busy = _add_tree_5_source_busy || _add_tree_5_sink_busy || _add_tree_5_busy_reg;
  reg _tmp_1816;
  reg _tmp_1817;
  reg _tmp_1818;
  reg _tmp_1819;
  reg _tmp_1820;
  reg _tmp_1821;
  reg _tmp_1822;
  reg _tmp_1823;
  reg _tmp_1824;
  reg _tmp_1825;
  assign _acc_1_source_stop = _acc_1_stream_oready && 1'd0;
  reg _tmp_1826;
  reg _tmp_1827;
  reg _tmp_1828;
  reg _tmp_1829;
  reg _tmp_1830;
  reg _tmp_1831;
  reg _tmp_1832;
  assign _acc_1_sink_start = _tmp_1832;
  reg _tmp_1833;
  reg _tmp_1834;
  reg _tmp_1835;
  reg _tmp_1836;
  reg _tmp_1837;
  reg _tmp_1838;
  reg _tmp_1839;
  assign _acc_1_sink_stop = _tmp_1839;
  reg _tmp_1840;
  reg _tmp_1841;
  reg _tmp_1842;
  reg _tmp_1843;
  reg _tmp_1844;
  reg _tmp_1845;
  reg _tmp_1846;
  assign _acc_1_sink_busy = _tmp_1846;
  reg _tmp_1847;
  assign _acc_1_busy = _acc_1_source_busy || _acc_1_sink_busy || _acc_1_busy_reg;
  reg _tmp_1848;
  reg _tmp_1849;
  reg _tmp_1850;
  assign _mul_rshift_round_clip_7_source_stop = _mul_rshift_round_clip_7_stream_oready && 1'd0;
  reg _tmp_1851;
  reg _tmp_1852;
  reg _tmp_1853;
  reg _tmp_1854;
  reg _tmp_1855;
  reg _tmp_1856;
  reg _tmp_1857;
  reg _tmp_1858;
  reg _tmp_1859;
  reg _tmp_1860;
  assign _mul_rshift_round_clip_7_sink_start = _tmp_1860;
  reg _tmp_1861;
  reg _tmp_1862;
  reg _tmp_1863;
  reg _tmp_1864;
  reg _tmp_1865;
  reg _tmp_1866;
  reg _tmp_1867;
  reg _tmp_1868;
  reg _tmp_1869;
  reg _tmp_1870;
  assign _mul_rshift_round_clip_7_sink_stop = _tmp_1870;
  reg _tmp_1871;
  reg _tmp_1872;
  reg _tmp_1873;
  reg _tmp_1874;
  reg _tmp_1875;
  reg _tmp_1876;
  reg _tmp_1877;
  reg _tmp_1878;
  reg _tmp_1879;
  reg _tmp_1880;
  assign _mul_rshift_round_clip_7_sink_busy = _tmp_1880;
  reg _tmp_1881;
  assign _mul_rshift_round_clip_7_busy = _mul_rshift_round_clip_7_source_busy || _mul_rshift_round_clip_7_sink_busy || _mul_rshift_round_clip_7_busy_reg;
  reg _tmp_1882;
  reg _tmp_1883;
  reg _tmp_1884;
  reg _tmp_1885;
  reg _tmp_1886;
  reg _tmp_1887;
  reg [1-1:0] __variable_wdata_951;
  assign stream_conv2d_4__reduce_reset_data = __variable_wdata_951;
  reg _tmp_1888;
  reg _tmp_1889;
  reg _tmp_1890;
  reg _tmp_1891;
  assign _stream_conv2d_4_source_stop = _stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_38_idle && _stream_conv2d_4_source_39_idle && _stream_conv2d_4_source_40_idle && _stream_conv2d_4_source_41_idle && _stream_conv2d_4_source_42_idle && _stream_conv2d_4_source_43_idle && _stream_conv2d_4_source_44_idle && _stream_conv2d_4_source_45_idle && _stream_conv2d_4_source_46_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3));
  localparam _tmp_1892 = 1;
  wire [_tmp_1892-1:0] _tmp_1893;
  assign _tmp_1893 = _stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_38_idle && _stream_conv2d_4_source_39_idle && _stream_conv2d_4_source_40_idle && _stream_conv2d_4_source_41_idle && _stream_conv2d_4_source_42_idle && _stream_conv2d_4_source_43_idle && _stream_conv2d_4_source_44_idle && _stream_conv2d_4_source_45_idle && _stream_conv2d_4_source_46_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3);
  reg [_tmp_1892-1:0] _tmp_1894;
  localparam _tmp_1895 = 1;
  wire [_tmp_1895-1:0] _tmp_1896;
  assign _tmp_1896 = _stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_38_idle && _stream_conv2d_4_source_39_idle && _stream_conv2d_4_source_40_idle && _stream_conv2d_4_source_41_idle && _stream_conv2d_4_source_42_idle && _stream_conv2d_4_source_43_idle && _stream_conv2d_4_source_44_idle && _stream_conv2d_4_source_45_idle && _stream_conv2d_4_source_46_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3);
  reg [_tmp_1895-1:0] _tmp_1897;
  reg _tmp_1898;
  reg _tmp_1899;
  reg _tmp_1900;
  reg _tmp_1901;
  reg _tmp_1902;
  reg _tmp_1903;
  reg _tmp_1904;
  reg _tmp_1905;
  reg _tmp_1906;
  reg _tmp_1907;
  reg _tmp_1908;
  reg _tmp_1909;
  reg _tmp_1910;
  reg _tmp_1911;
  reg _tmp_1912;
  reg _tmp_1913;
  reg _tmp_1914;
  reg _tmp_1915;
  reg _tmp_1916;
  reg _tmp_1917;
  reg _tmp_1918;
  reg _tmp_1919;
  reg _tmp_1920;
  reg _tmp_1921;
  reg _tmp_1922;
  reg _tmp_1923;
  reg _tmp_1924;
  reg _tmp_1925;
  reg _tmp_1926;
  reg _tmp_1927;
  reg _tmp_1928;
  reg _tmp_1929;
  reg _tmp_1930;
  reg _tmp_1931;
  reg _tmp_1932;
  reg _tmp_1933;
  assign _stream_conv2d_4_sink_start = _tmp_1933;
  reg _tmp_1934;
  reg _tmp_1935;
  reg _tmp_1936;
  reg _tmp_1937;
  reg _tmp_1938;
  reg _tmp_1939;
  reg _tmp_1940;
  reg _tmp_1941;
  reg _tmp_1942;
  reg _tmp_1943;
  reg _tmp_1944;
  reg _tmp_1945;
  reg _tmp_1946;
  reg _tmp_1947;
  reg _tmp_1948;
  reg _tmp_1949;
  reg _tmp_1950;
  reg _tmp_1951;
  reg _tmp_1952;
  reg _tmp_1953;
  reg _tmp_1954;
  reg _tmp_1955;
  reg _tmp_1956;
  reg _tmp_1957;
  reg _tmp_1958;
  reg _tmp_1959;
  reg _tmp_1960;
  reg _tmp_1961;
  reg _tmp_1962;
  reg _tmp_1963;
  reg _tmp_1964;
  reg _tmp_1965;
  reg _tmp_1966;
  reg _tmp_1967;
  reg _tmp_1968;
  reg _tmp_1969;
  assign _stream_conv2d_4_sink_stop = _tmp_1969;
  reg _tmp_1970;
  reg _tmp_1971;
  reg _tmp_1972;
  reg _tmp_1973;
  reg _tmp_1974;
  reg _tmp_1975;
  reg _tmp_1976;
  reg _tmp_1977;
  reg _tmp_1978;
  reg _tmp_1979;
  reg _tmp_1980;
  reg _tmp_1981;
  reg _tmp_1982;
  reg _tmp_1983;
  reg _tmp_1984;
  reg _tmp_1985;
  reg _tmp_1986;
  reg _tmp_1987;
  reg _tmp_1988;
  reg _tmp_1989;
  reg _tmp_1990;
  reg _tmp_1991;
  reg _tmp_1992;
  reg _tmp_1993;
  reg _tmp_1994;
  reg _tmp_1995;
  reg _tmp_1996;
  reg _tmp_1997;
  reg _tmp_1998;
  reg _tmp_1999;
  reg _tmp_2000;
  reg _tmp_2001;
  reg _tmp_2002;
  reg _tmp_2003;
  reg _tmp_2004;
  reg _tmp_2005;
  assign _stream_conv2d_4_sink_busy = _tmp_2005;
  reg _tmp_2006;
  assign _stream_conv2d_4_busy = _stream_conv2d_4_source_busy || _stream_conv2d_4_sink_busy || _stream_conv2d_4_busy_reg;
  wire conv2d_4_dma_out_mask_0;
  assign conv2d_4_dma_out_mask_0 = conv2d_4_out_row_count + 0 >= cparam_conv2d_4_out_num_row;
  wire [32-1:0] mask_addr_shifted_2007;
  assign mask_addr_shifted_2007 = conv2d_4_objaddr + (conv2d_4_out_base_offset + cparam_conv2d_4_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2008;
  assign mask_addr_masked_2008 = mask_addr_shifted_2007 << 2;
  reg [32-1:0] _maxi_write_req_fsm;
  localparam _maxi_write_req_fsm_init = 0;
  reg [33-1:0] _maxi_write_cur_global_size;
  reg _maxi_write_cont;
  wire [8-1:0] pack_write_req_op_sel_2009;
  wire [32-1:0] pack_write_req_local_addr_2010;
  wire [32-1:0] pack_write_req_local_stride_2011;
  wire [33-1:0] pack_write_req_size_2012;
  wire [32-1:0] pack_write_req_local_blocksize_2013;
  assign pack_write_req_op_sel_2009 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_2010 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_2011 = _maxi_write_local_stride;
  assign pack_write_req_size_2012 = _maxi_write_local_size;
  assign pack_write_req_local_blocksize_2013 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_2014;
  assign pack_write_req_packed_2014 = { pack_write_req_op_sel_2009, pack_write_req_local_addr_2010, pack_write_req_local_stride_2011, pack_write_req_size_2012, pack_write_req_local_blocksize_2013 };
  localparam _tmp_2015 = 1;
  wire [_tmp_2015-1:0] _tmp_2016;
  assign _tmp_2016 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_2015-1:0] __tmp_2016_1;
  wire [32-1:0] mask_addr_shifted_2017;
  assign mask_addr_shifted_2017 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_2018;
  assign mask_addr_masked_2018 = mask_addr_shifted_2017 << 2;
  wire [32-1:0] mask_addr_shifted_2019;
  assign mask_addr_shifted_2019 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_2020;
  assign mask_addr_masked_2020 = mask_addr_shifted_2019 << 2;
  wire [32-1:0] mask_addr_shifted_2021;
  assign mask_addr_shifted_2021 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_2022;
  assign mask_addr_masked_2022 = mask_addr_shifted_2021 << 2;
  wire [32-1:0] mask_addr_shifted_2023;
  assign mask_addr_shifted_2023 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_2024;
  assign mask_addr_masked_2024 = mask_addr_shifted_2023 << 2;
  wire [32-1:0] mask_addr_shifted_2025;
  assign mask_addr_shifted_2025 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_2026;
  assign mask_addr_masked_2026 = mask_addr_shifted_2025 << 2;
  wire [32-1:0] mask_addr_shifted_2027;
  assign mask_addr_shifted_2027 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_2028;
  assign mask_addr_masked_2028 = mask_addr_shifted_2027 << 2;
  wire [8-1:0] pack_write_req_op_sel_2029;
  wire [32-1:0] pack_write_req_local_addr_2030;
  wire [32-1:0] pack_write_req_local_stride_2031;
  wire [33-1:0] pack_write_req_size_2032;
  wire [32-1:0] pack_write_req_local_blocksize_2033;
  assign pack_write_req_op_sel_2029 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_2030 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_2031 = _maxi_write_local_stride;
  assign pack_write_req_size_2032 = _maxi_write_cur_global_size;
  assign pack_write_req_local_blocksize_2033 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_2034;
  assign pack_write_req_packed_2034 = { pack_write_req_op_sel_2029, pack_write_req_local_addr_2030, pack_write_req_local_stride_2031, pack_write_req_size_2032, pack_write_req_local_blocksize_2033 };
  assign _maxi_write_req_fifo_wdata = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? pack_write_req_packed_2034 : 
                                      ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? pack_write_req_packed_2014 : 'hx;
  assign _maxi_write_req_fifo_enq = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? (_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && !_maxi_write_req_fifo_almost_full : 
                                    ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? (_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full && !_maxi_write_req_fifo_almost_full : 0;
  localparam _tmp_2035 = 1;
  wire [_tmp_2035-1:0] _tmp_2036;
  assign _tmp_2036 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_2035-1:0] __tmp_2036_1;
  reg _maxi_waddr_cond_0_1;
  reg [32-1:0] _maxi_write_data_fsm;
  localparam _maxi_write_data_fsm_init = 0;
  reg [32-1:0] read_burst_fsm_33;
  localparam read_burst_fsm_33_init = 0;
  reg [7-1:0] read_burst_addr_2037;
  reg [7-1:0] read_burst_stride_2038;
  reg [33-1:0] read_burst_length_2039;
  reg read_burst_rvalid_2040;
  reg read_burst_rlast_2041;
  assign ram_w32_l128_id20_1_addr = ((read_burst_fsm_33 == 1) && (!read_burst_rvalid_2040 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_2037 : 'hx;
  assign ram_w32_l128_id20_1_enable = ((read_burst_fsm_33 == 1) && (!read_burst_rvalid_2040 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_2042 = 1;
  wire [_tmp_2042-1:0] _tmp_2043;
  assign _tmp_2043 = (read_burst_fsm_33 == 1) && (!read_burst_rvalid_2040 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_2042-1:0] __tmp_2043_1;
  wire [32-1:0] read_burst_rdata_2044;
  assign read_burst_rdata_2044 = ram_w32_l128_id20_1_rdata;
  reg _maxi_wdata_cond_0_1;
  wire conv2d_4_update_filter;
  assign conv2d_4_update_filter = (cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) || (cparam_conv2d_4_data_stationary == 1) && !cparam_conv2d_4_keep_filter;
  wire conv2d_4_update_act;
  assign conv2d_4_update_act = (cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) || (cparam_conv2d_4_data_stationary == 0);
  wire conv2d_4_mux_next_dma_flag_0;
  assign conv2d_4_mux_next_dma_flag_0 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 1'd0;
  wire conv2d_4_mux_next_dma_flag_1;
  assign conv2d_4_mux_next_dma_flag_1 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 1'd0;
  wire conv2d_4_mux_next_dma_flag_2;
  assign conv2d_4_mux_next_dma_flag_2 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] max_pool_serial_6_objaddr;
  reg [32-1:0] max_pool_serial_6_arg_objaddr_0;
  reg [32-1:0] control_max_pool_serial_6;
  localparam control_max_pool_serial_6_init = 0;
  reg _control_max_pool_serial_6_called;
  wire signed [32-1:0] max_pool_serial_6_act_base_offset;
  reg signed [32-1:0] max_pool_serial_6_act_base_offset_row;
  reg signed [32-1:0] max_pool_serial_6_act_base_offset_bat;
  assign max_pool_serial_6_act_base_offset = max_pool_serial_6_act_base_offset_row + max_pool_serial_6_act_base_offset_bat;
  wire signed [32-1:0] max_pool_serial_6_out_base_offset;
  reg signed [32-1:0] max_pool_serial_6_out_base_offset_row;
  reg signed [32-1:0] max_pool_serial_6_out_base_offset_bat;
  assign max_pool_serial_6_out_base_offset = max_pool_serial_6_out_base_offset_row + max_pool_serial_6_out_base_offset_bat;
  reg [32-1:0] max_pool_serial_6_col_count;
  reg [32-1:0] max_pool_serial_6_row_count;
  reg [32-1:0] max_pool_serial_6_bat_count;
  reg [32-1:0] max_pool_serial_6_prev_row_count;
  reg [32-1:0] max_pool_serial_6_prev_bat_count;
  reg [32-1:0] max_pool_serial_6_stream_act_local;
  reg [32-1:0] max_pool_serial_6_stream_out_local;
  reg max_pool_serial_6_act_page;
  reg [32-1:0] max_pool_serial_6_act_page_comp_offset;
  reg [32-1:0] max_pool_serial_6_act_page_dma_offset;
  reg max_pool_serial_6_out_page;
  reg [32-1:0] max_pool_serial_6_out_page_comp_offset;
  reg [32-1:0] max_pool_serial_6_out_page_dma_offset;
  reg max_pool_serial_6_skip_read_act;
  reg max_pool_serial_6_skip_comp;
  reg max_pool_serial_6_skip_write_out;
  reg [32-1:0] max_pool_serial_6_comp_count;
  reg [32-1:0] max_pool_serial_6_out_count;
  wire max_pool_serial_6_dma_pad_mask_0;
  assign max_pool_serial_6_dma_pad_mask_0 = (max_pool_serial_6_row_count + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_dma_pad_mask_1;
  assign max_pool_serial_6_dma_pad_mask_1 = (max_pool_serial_6_row_count + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire [32-1:0] mask_addr_shifted_2045;
  assign mask_addr_shifted_2045 = max_pool_serial_6_arg_objaddr_0 + (max_pool_serial_6_act_base_offset + cparam_max_pool_serial_6_act_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2046;
  assign mask_addr_masked_2046 = mask_addr_shifted_2045 << 2;
  reg [32-1:0] write_burst_fsm_34;
  localparam write_burst_fsm_34_init = 0;
  reg [14-1:0] write_burst_addr_2047;
  reg [14-1:0] write_burst_stride_2048;
  reg [33-1:0] write_burst_length_2049;
  reg write_burst_done_2050;
  wire [32-1:0] mask_addr_shifted_2051;
  assign mask_addr_shifted_2051 = max_pool_serial_6_arg_objaddr_0 + (max_pool_serial_6_act_base_offset + cparam_max_pool_serial_6_act_offset_values_1) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2052;
  assign mask_addr_masked_2052 = mask_addr_shifted_2051 << 2;
  reg [32-1:0] max_pool_serial_6_comp_fsm;
  localparam max_pool_serial_6_comp_fsm_init = 0;
  reg [32-1:0] max_pool_serial_6_act_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_6_out_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_6_row_count_buf;
  wire max_pool_serial_6_stream_pad_mask_0_0;
  assign max_pool_serial_6_stream_pad_mask_0_0 = (max_pool_serial_6_col_count + 0 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 0 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_0_1;
  assign max_pool_serial_6_stream_pad_mask_0_1 = (max_pool_serial_6_col_count + 1 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 1 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_1_0;
  assign max_pool_serial_6_stream_pad_mask_1_0 = (max_pool_serial_6_col_count + 0 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 0 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_1_1;
  assign max_pool_serial_6_stream_pad_mask_1_1 = (max_pool_serial_6_col_count + 1 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 1 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  reg [4-1:0] max_pool_serial_6_stream_pad_masks;
  wire [3-1:0] stream_max_pool_serial_6_parameter_0_data;
  wire [32-1:0] stream_max_pool_serial_6_source_1_data;
  wire [4-1:0] stream_max_pool_serial_6_parameter_2_data;
  wire [1-1:0] stream_max_pool_serial_6__reduce_reset_data;
  reg __stream_max_pool_serial_6_stream_ivalid_1;
  reg __stream_max_pool_serial_6_stream_ivalid_2;
  reg __stream_max_pool_serial_6_stream_ivalid_3;
  reg __stream_max_pool_serial_6_stream_ivalid_4;
  reg __stream_max_pool_serial_6_stream_ivalid_5;
  reg [32-1:0] _counter_data_2421;
  reg [32-1:0] _counter_count_2421;
  wire _counter_reset_cond_2421;
  assign _counter_reset_cond_2421 = stream_max_pool_serial_6__reduce_reset_data;
  wire [32-1:0] _counter_current_count_2421;
  assign _counter_current_count_2421 = (_counter_reset_cond_2421)? 1'sd0 : _counter_count_2421;
  wire [16-1:0] _slice_data_2427;
  assign _slice_data_2427 = stream_max_pool_serial_6_source_1_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2428;
  assign _reinterpretcast_src_2428 = _slice_data_2427;
  wire signed [16-1:0] _reinterpretcast_data_2428;
  assign _reinterpretcast_data_2428 = _reinterpretcast_src_2428;
  wire [16-1:0] _slice_data_2431;
  assign _slice_data_2431 = stream_max_pool_serial_6_source_1_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2432;
  assign _reinterpretcast_src_2432 = _slice_data_2431;
  wire signed [16-1:0] _reinterpretcast_data_2432;
  assign _reinterpretcast_data_2432 = _reinterpretcast_src_2432;
  reg [4-1:0] __delay_data_3108__variable_2419;
  reg signed [16-1:0] __delay_data_3109_reinterpretcast_2428;
  reg [1-1:0] __delay_data_3111__variable_2420;
  reg [3-1:0] __delay_data_3114__variable_2417;
  reg signed [16-1:0] __delay_data_3117_reinterpretcast_2432;
  reg [1-1:0] _pointer_data_2424;
  reg signed [16-1:0] __delay_data_3110__delay_3109_reinterpretcast_2428;
  reg [1-1:0] __delay_data_3112__delay_3111__variable_2420;
  reg [3-1:0] __delay_data_3115__delay_3114__variable_2417;
  reg signed [16-1:0] __delay_data_3118__delay_3117_reinterpretcast_2432;
  reg signed [17-1:0] _cond_data_2434;
  reg signed [17-1:0] _cond_data_2439;
  reg [1-1:0] __delay_data_3113__delay_3112__delay_3111__variable_2420;
  reg [3-1:0] __delay_data_3116__delay_3115__delay_3114__variable_2417;
  reg [1-1:0] __variable_wdata_934;
  assign _reduce_max_44__reduce_reset_data = __variable_wdata_934;
  reg signed [16-1:0] __variable_wdata_932;
  assign _reduce_max_44_x_data = __variable_wdata_932;
  reg [32-1:0] __variable_wdata_933;
  assign _reduce_max_44_size_data = __variable_wdata_933;
  assign __reduce_max_44_is_root = ((_stream_max_pool_serial_6_busy)? 0 : 1) && 1;
  assign __reduce_max_44_stream_oready = ((_stream_max_pool_serial_6_busy)? _stream_max_pool_serial_6_stream_oready : 1) && __reduce_max_44_stream_internal_oready;
  reg [1-1:0] __variable_wdata_941;
  assign _reduce_max_45__reduce_reset_data = __variable_wdata_941;
  reg signed [16-1:0] __variable_wdata_939;
  assign _reduce_max_45_x_data = __variable_wdata_939;
  reg [32-1:0] __variable_wdata_940;
  assign _reduce_max_45_size_data = __variable_wdata_940;
  assign __reduce_max_45_is_root = ((_stream_max_pool_serial_6_busy)? 0 : 1) && 1;
  assign __reduce_max_45_stream_oready = ((_stream_max_pool_serial_6_busy)? _stream_max_pool_serial_6_stream_oready : 1) && __reduce_max_45_stream_internal_oready;
  assign _stream_max_pool_serial_6_stream_internal_oready = ((_stream_max_pool_serial_6_busy)? __reduce_max_45_stream_internal_oready : 1) && (((_stream_max_pool_serial_6_busy)? __reduce_max_44_stream_internal_oready : 1) && 1);
  wire signed [16-1:0] __substreamoutput_data_2436;
  assign __substreamoutput_data_2436 = _reduce_max_44_data_data;
  wire [1-1:0] __substreamoutput_data_2437;
  assign __substreamoutput_data_2437 = _reduce_max_44_valid_data;
  wire signed [16-1:0] _reinterpretcast_src_2438;
  assign _reinterpretcast_src_2438 = __substreamoutput_data_2436;
  wire signed [16-1:0] _reinterpretcast_data_2438;
  assign _reinterpretcast_data_2438 = _reinterpretcast_src_2438;
  wire signed [16-1:0] __substreamoutput_data_2441;
  assign __substreamoutput_data_2441 = _reduce_max_45_data_data;
  wire signed [16-1:0] _reinterpretcast_src_2443;
  assign _reinterpretcast_src_2443 = __substreamoutput_data_2441;
  wire signed [16-1:0] _reinterpretcast_data_2443;
  assign _reinterpretcast_data_2443 = _reinterpretcast_src_2443;
  wire [32-1:0] _cat_data_2444;
  assign _cat_data_2444 = { _reinterpretcast_data_2443, _reinterpretcast_data_2438 };
  wire [1-1:0] stream_max_pool_serial_6_sink_7_data;
  assign stream_max_pool_serial_6_sink_7_data = __substreamoutput_data_2437;
  wire [32-1:0] stream_max_pool_serial_6_sink_6_data;
  assign stream_max_pool_serial_6_sink_6_data = _cat_data_2444;
  wire _set_flag_2053;
  assign _set_flag_2053 = max_pool_serial_6_comp_fsm == 4;
  reg [3-1:0] __variable_wdata_2417;
  assign stream_max_pool_serial_6_parameter_0_data = __variable_wdata_2417;
  wire _set_flag_2054;
  assign _set_flag_2054 = max_pool_serial_6_comp_fsm == 4;
  reg [4-1:0] __variable_wdata_2419;
  assign stream_max_pool_serial_6_parameter_2_data = __variable_wdata_2419;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_3;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_3;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3;
  wire _set_flag_2055;
  assign _set_flag_2055 = max_pool_serial_6_comp_fsm == 4;
  localparam _tmp_2056 = 1;
  wire [_tmp_2056-1:0] _tmp_2057;
  assign _tmp_2057 = _stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1);
  reg [_tmp_2056-1:0] __tmp_2057_1;
  assign _stream_max_pool_serial_6_source_1_source_ram_rdata = (_stream_max_pool_serial_6_source_1_source_sel == 1)? ram_w32_l16384_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_2418;
  assign stream_max_pool_serial_6_source_1_data = __variable_wdata_2418;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_pat_fsm_0;
  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_max_pool_serial_6_source_1_source_pat_all_offset;
  assign _stream_max_pool_serial_6_source_1_source_pat_all_offset = _stream_max_pool_serial_6_source_1_source_offset_buf + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3;
  wire _set_flag_2058;
  assign _set_flag_2058 = max_pool_serial_6_comp_fsm == 4;
  reg _tmp_2059;
  reg _tmp_2060;
  reg _tmp_2061;
  reg _tmp_2062;
  reg _tmp_2063;
  reg _tmp_2064;
  reg _tmp_2065;
  localparam _tmp_2066 = 33;
  wire [_tmp_2066-1:0] _tmp_2067;
  assign _tmp_2067 = max_pool_serial_6_stream_out_local + max_pool_serial_6_out_page_comp_offset_buf;
  reg [_tmp_2066-1:0] _tmp_2068;
  reg [_tmp_2066-1:0] _tmp_2069;
  reg [_tmp_2066-1:0] _tmp_2070;
  reg [_tmp_2066-1:0] _tmp_2071;
  reg [_tmp_2066-1:0] _tmp_2072;
  reg [_tmp_2066-1:0] _tmp_2073;
  reg [_tmp_2066-1:0] _tmp_2074;
  reg [6-1:0] _tmp_2075;
  reg [6-1:0] _tmp_2076;
  reg [6-1:0] _tmp_2077;
  reg [6-1:0] _tmp_2078;
  reg [6-1:0] _tmp_2079;
  reg [6-1:0] _tmp_2080;
  reg [6-1:0] _tmp_2081;
  assign ram_w32_l8192_id0_0_wdata = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? _stream_max_pool_serial_6_sink_6_sink_wdata : 'hx;
  assign ram_w32_l8192_id0_0_wenable = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? 1'd1 : 0;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_fsm_1;
  localparam _stream_max_pool_serial_6_sink_6_sink_fsm_1_init = 0;
  wire _set_flag_2082;
  assign _set_flag_2082 = max_pool_serial_6_comp_fsm == 5;
  assign _stream_max_pool_serial_6_run_flag = (_set_flag_2082)? 1 : 0;
  reg _tmp_2083;
  reg _tmp_2084;
  reg _tmp_2085;
  reg _tmp_2086;
  reg _tmp_2087;
  reg _tmp_2088;
  reg _tmp_2089;
  reg _tmp_2090;
  reg _tmp_2091;
  reg _tmp_2092;
  assign __reduce_max_44_source_stop = __reduce_max_44_stream_oready && 1'd0;
  reg _tmp_2093;
  reg _tmp_2094;
  reg _tmp_2095;
  assign __reduce_max_44_sink_start = _tmp_2095;
  reg _tmp_2096;
  reg _tmp_2097;
  reg _tmp_2098;
  assign __reduce_max_44_sink_stop = _tmp_2098;
  reg _tmp_2099;
  reg _tmp_2100;
  reg _tmp_2101;
  assign __reduce_max_44_sink_busy = _tmp_2101;
  reg _tmp_2102;
  assign __reduce_max_44_busy = __reduce_max_44_source_busy || __reduce_max_44_sink_busy || __reduce_max_44_busy_reg;
  reg _tmp_2103;
  reg _tmp_2104;
  reg _tmp_2105;
  reg _tmp_2106;
  reg _tmp_2107;
  reg _tmp_2108;
  reg _tmp_2109;
  reg _tmp_2110;
  reg _tmp_2111;
  reg _tmp_2112;
  assign __reduce_max_45_source_stop = __reduce_max_45_stream_oready && 1'd0;
  reg _tmp_2113;
  reg _tmp_2114;
  reg _tmp_2115;
  assign __reduce_max_45_sink_start = _tmp_2115;
  reg _tmp_2116;
  reg _tmp_2117;
  reg _tmp_2118;
  assign __reduce_max_45_sink_stop = _tmp_2118;
  reg _tmp_2119;
  reg _tmp_2120;
  reg _tmp_2121;
  assign __reduce_max_45_sink_busy = _tmp_2121;
  reg _tmp_2122;
  assign __reduce_max_45_busy = __reduce_max_45_source_busy || __reduce_max_45_sink_busy || __reduce_max_45_busy_reg;
  reg _tmp_2123;
  reg _tmp_2124;
  reg _tmp_2125;
  reg _tmp_2126;
  reg _tmp_2127;
  reg _tmp_2128;
  reg [1-1:0] __variable_wdata_2420;
  assign stream_max_pool_serial_6__reduce_reset_data = __variable_wdata_2420;
  reg _tmp_2129;
  reg _tmp_2130;
  reg _tmp_2131;
  reg _tmp_2132;
  assign _stream_max_pool_serial_6_source_stop = _stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3));
  localparam _tmp_2133 = 1;
  wire [_tmp_2133-1:0] _tmp_2134;
  assign _tmp_2134 = _stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3);
  reg [_tmp_2133-1:0] _tmp_2135;
  localparam _tmp_2136 = 1;
  wire [_tmp_2136-1:0] _tmp_2137;
  assign _tmp_2137 = _stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3);
  reg [_tmp_2136-1:0] _tmp_2138;
  reg _tmp_2139;
  reg _tmp_2140;
  reg _tmp_2141;
  reg _tmp_2142;
  reg _tmp_2143;
  reg _tmp_2144;
  reg _tmp_2145;
  assign _stream_max_pool_serial_6_sink_start = _tmp_2145;
  reg _tmp_2146;
  reg _tmp_2147;
  reg _tmp_2148;
  reg _tmp_2149;
  reg _tmp_2150;
  reg _tmp_2151;
  reg _tmp_2152;
  assign _stream_max_pool_serial_6_sink_stop = _tmp_2152;
  reg _tmp_2153;
  reg _tmp_2154;
  reg _tmp_2155;
  reg _tmp_2156;
  reg _tmp_2157;
  reg _tmp_2158;
  reg _tmp_2159;
  assign _stream_max_pool_serial_6_sink_busy = _tmp_2159;
  reg _tmp_2160;
  assign _stream_max_pool_serial_6_busy = _stream_max_pool_serial_6_source_busy || _stream_max_pool_serial_6_sink_busy || _stream_max_pool_serial_6_busy_reg;
  wire [32-1:0] mask_addr_shifted_2161;
  assign mask_addr_shifted_2161 = max_pool_serial_6_objaddr + max_pool_serial_6_out_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2162;
  assign mask_addr_masked_2162 = mask_addr_shifted_2161 << 2;
  reg [32-1:0] read_burst_fsm_35;
  localparam read_burst_fsm_35_init = 0;
  reg [13-1:0] read_burst_addr_2163;
  reg [13-1:0] read_burst_stride_2164;
  reg [33-1:0] read_burst_length_2165;
  reg read_burst_rvalid_2166;
  reg read_burst_rlast_2167;
  localparam _tmp_2168 = 1;
  wire [_tmp_2168-1:0] _tmp_2169;
  assign _tmp_2169 = (read_burst_fsm_35 == 1) && (!read_burst_rvalid_2166 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_2168-1:0] __tmp_2169_1;
  wire [32-1:0] read_burst_rdata_2170;
  assign read_burst_rdata_2170 = ram_w32_l8192_id0_1_rdata;
  reg _maxi_wdata_cond_1_1;
  reg [32-1:0] matmul_16_objaddr;
  reg [32-1:0] matmul_16_arg_objaddr_0;
  reg [32-1:0] matmul_16_arg_objaddr_1;
  reg [32-1:0] matmul_16_arg_objaddr_2;
  reg [32-1:0] matmul_16_arg_objaddr_3;
  reg [32-1:0] control_matmul_16;
  localparam control_matmul_16_init = 0;
  reg _control_matmul_16_called;
  wire signed [32-1:0] matmul_16_act_base_offset;
  reg signed [32-1:0] matmul_16_act_base_offset_row;
  reg signed [32-1:0] matmul_16_act_base_offset_bat;
  assign matmul_16_act_base_offset = matmul_16_act_base_offset_row + matmul_16_act_base_offset_bat;
  reg signed [32-1:0] matmul_16_filter_base_offset;
  reg [32-1:0] matmul_16_next_stream_num_ops;
  wire signed [32-1:0] matmul_16_out_base_offset;
  reg signed [32-1:0] matmul_16_out_base_offset_val;
  reg signed [32-1:0] matmul_16_out_base_offset_col;
  reg signed [32-1:0] matmul_16_out_base_offset_row;
  reg signed [32-1:0] matmul_16_out_base_offset_bat;
  reg signed [32-1:0] matmul_16_out_base_offset_och;
  assign matmul_16_out_base_offset = matmul_16_out_base_offset_val + matmul_16_out_base_offset_col + matmul_16_out_base_offset_row + matmul_16_out_base_offset_bat + matmul_16_out_base_offset_och;
  reg matmul_16_dma_flag_0;
  reg [32-1:0] matmul_16_sync_comp_count;
  reg [32-1:0] matmul_16_sync_out_count;
  reg [32-1:0] matmul_16_write_count;
  reg [32-1:0] matmul_16_next_out_write_size;
  reg [32-1:0] matmul_16_col_count;
  reg [32-1:0] matmul_16_row_count;
  reg [32-1:0] matmul_16_bat_count;
  reg [32-1:0] matmul_16_och_count;
  reg [1-1:0] matmul_16_col_select;
  reg [1-1:0] matmul_16_row_select;
  reg [32-1:0] matmul_16_out_col_count;
  reg [32-1:0] matmul_16_out_row_count;
  reg [32-1:0] matmul_16_out_ram_select;
  reg [32-1:0] matmul_16_prev_col_count;
  reg [32-1:0] matmul_16_prev_row_count;
  reg [32-1:0] matmul_16_prev_bat_count;
  reg [32-1:0] matmul_16_prev_och_count;
  reg [1-1:0] matmul_16_prev_row_select;
  reg [32-1:0] matmul_16_stream_act_local_0;
  reg [32-1:0] matmul_16_stream_out_local_val;
  reg [32-1:0] matmul_16_stream_out_local_col;
  wire [32-1:0] matmul_16_stream_out_local;
  assign matmul_16_stream_out_local = matmul_16_stream_out_local_val + matmul_16_stream_out_local_col;
  reg [32-1:0] matmul_16_act_page_comp_offset_0;
  reg [32-1:0] matmul_16_act_page_dma_offset_0;
  reg [32-1:0] matmul_16_filter_page_comp_offset;
  reg [32-1:0] matmul_16_filter_page_dma_offset;
  reg matmul_16_out_page;
  reg [32-1:0] matmul_16_out_page_comp_offset;
  reg [32-1:0] matmul_16_out_page_dma_offset;
  reg [32-1:0] matmul_16_out_laddr_offset;
  reg matmul_16_skip_read_filter;
  reg matmul_16_skip_read_act;
  reg matmul_16_skip_comp;
  reg matmul_16_skip_write_out;
  wire [32-1:0] mask_addr_shifted_2171;
  assign mask_addr_shifted_2171 = matmul_16_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2172;
  assign mask_addr_masked_2172 = mask_addr_shifted_2171 << 2;
  reg [32-1:0] write_burst_fsm_36;
  localparam write_burst_fsm_36_init = 0;
  reg [8-1:0] write_burst_addr_2173;
  reg [8-1:0] write_burst_stride_2174;
  reg [33-1:0] write_burst_length_2175;
  reg write_burst_done_2176;
  assign ram_w32_l256_id0_1_addr = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_2173 : 'hx;
  assign ram_w32_l256_id0_1_wdata = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l256_id0_1_wenable = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l256_id0_1_enable = ((write_burst_fsm_36 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_2177;
  assign mask_addr_shifted_2177 = matmul_16_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2178;
  assign mask_addr_masked_2178 = mask_addr_shifted_2177 << 2;
  reg [32-1:0] write_burst_fsm_37;
  localparam write_burst_fsm_37_init = 0;
  reg [8-1:0] write_burst_addr_2179;
  reg [8-1:0] write_burst_stride_2180;
  reg [33-1:0] write_burst_length_2181;
  reg write_burst_done_2182;
  assign ram_w32_l256_id1_1_addr = ((write_burst_fsm_37 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_2179 : 'hx;
  assign ram_w32_l256_id1_1_wdata = ((write_burst_fsm_37 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l256_id1_1_wenable = ((write_burst_fsm_37 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l256_id1_1_enable = ((write_burst_fsm_37 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_2183;
  assign mask_addr_shifted_2183 = matmul_16_arg_objaddr_1 + matmul_16_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2184;
  assign mask_addr_masked_2184 = mask_addr_shifted_2183 << 2;
  wire write_burst_block_ram_wvalid_2185;
  wire write_burst_block_ram_wquit_2186;
  reg [32-1:0] write_burst_fsm_38;
  localparam write_burst_fsm_38_init = 0;
  reg [14-1:0] write_burst_addr_2187;
  reg [14-1:0] write_burst_stride_2188;
  reg [33-1:0] write_burst_length_2189;
  reg write_burst_done_2190;
  assign ram_w32_l16384_id0_1_addr = ((write_burst_fsm_38 == 1) && write_burst_block_ram_wvalid_2185)? write_burst_addr_2187 : 
                                     ((write_burst_fsm_34 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_2047 : 'hx;
  assign ram_w32_l16384_id0_1_wdata = ((write_burst_fsm_38 == 1) && write_burst_block_ram_wvalid_2185)? _maxi_rdata_sb_0 : 
                                      ((write_burst_fsm_34 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l16384_id0_1_wenable = ((write_burst_fsm_38 == 1) && write_burst_block_ram_wvalid_2185)? 1'd1 : 
                                        ((write_burst_fsm_34 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l16384_id0_1_enable = ((write_burst_fsm_38 == 1) && write_burst_block_ram_wvalid_2185)? 1'd1 : 
                                       ((write_burst_fsm_34 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_2191;
  wire write_burst_block_ram_wquit_2192;
  reg [32-1:0] write_burst_fsm_39;
  localparam write_burst_fsm_39_init = 0;
  reg [14-1:0] write_burst_addr_2193;
  reg [14-1:0] write_burst_stride_2194;
  reg [33-1:0] write_burst_length_2195;
  reg write_burst_done_2196;
  assign ram_w32_l16384_id1_1_addr = ((write_burst_fsm_39 == 1) && write_burst_block_ram_wvalid_2191)? write_burst_addr_2193 : 'hx;
  assign ram_w32_l16384_id1_1_wdata = ((write_burst_fsm_39 == 1) && write_burst_block_ram_wvalid_2191)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l16384_id1_1_wenable = ((write_burst_fsm_39 == 1) && write_burst_block_ram_wvalid_2191)? 1'd1 : 0;
  assign ram_w32_l16384_id1_1_enable = ((write_burst_fsm_39 == 1) && write_burst_block_ram_wvalid_2191)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_40;
  localparam write_burst_block_fsm_40_init = 0;
  reg [33-1:0] write_burst_block_length_2197;
  reg [32-1:0] write_burst_block_blocksize_2198;
  reg write_burst_block_done_2199;
  reg [32-1:0] write_burst_block_count_2200;
  assign write_burst_block_ram_wvalid_2185 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_40 == 1);
  assign write_burst_block_ram_wquit_2186 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_2197 <= 1);
  assign write_burst_block_ram_wvalid_2191 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_40 == 2);
  assign write_burst_block_ram_wquit_2192 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_2197 <= 1);
  wire [32-1:0] matmul_16_mux_act_gaddr_0;
  assign matmul_16_mux_act_gaddr_0 = (matmul_16_row_select == 0)? matmul_16_arg_objaddr_0 + (matmul_16_act_base_offset + cparam_matmul_16_act_offset_values_0) : 1'd0;
  wire matmul_16_dma_pad_mask_0;
  assign matmul_16_dma_pad_mask_0 = (matmul_16_row_count + 0 < cparam_matmul_16_pad_row_top) || (matmul_16_row_count + 0 >= cparam_matmul_16_act_num_row + cparam_matmul_16_pad_row_top);
  wire matmul_16_mux_dma_pad_mask_0;
  assign matmul_16_mux_dma_pad_mask_0 = (matmul_16_row_select == 0)? matmul_16_dma_pad_mask_0 : 1'd0;
  wire matmul_16_mux_dma_flag_0;
  assign matmul_16_mux_dma_flag_0 = (matmul_16_prev_row_select == 0)? matmul_16_dma_flag_0 : 1'd0;
  wire [32-1:0] mask_addr_shifted_2201;
  assign mask_addr_shifted_2201 = matmul_16_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2202;
  assign mask_addr_masked_2202 = mask_addr_shifted_2201 << 2;
  assign _maxi_read_req_fifo_deq = ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 11)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) && !_maxi_read_req_fifo_empty)? 1 : 0;
  reg [32-1:0] write_burst_fsm_41;
  localparam write_burst_fsm_41_init = 0;
  reg [13-1:0] write_burst_addr_2203;
  reg [13-1:0] write_burst_stride_2204;
  reg [33-1:0] write_burst_length_2205;
  reg write_burst_done_2206;
  assign ram_w32_l8192_id0_1_addr = ((write_burst_fsm_41 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_2203 : 
                                    ((read_burst_fsm_35 == 1) && (!read_burst_rvalid_2166 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_2163 : 'hx;
  assign ram_w32_l8192_id0_1_wdata = ((write_burst_fsm_41 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l8192_id0_1_wenable = ((write_burst_fsm_41 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l8192_id0_1_enable = ((write_burst_fsm_41 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                      ((read_burst_fsm_35 == 1) && (!read_burst_rvalid_2166 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  assign _maxi_rready_sb_0 = (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2);
  reg [32-1:0] matmul_16_comp_fsm;
  localparam matmul_16_comp_fsm_init = 0;
  reg [32-1:0] matmul_16_filter_page_comp_offset_buf;
  reg [32-1:0] matmul_16_act_page_comp_offset_buf_0;
  reg [32-1:0] matmul_16_out_page_comp_offset_buf;
  reg [32-1:0] matmul_16_row_count_buf;
  reg [1-1:0] matmul_16_row_select_buf;
  reg [32-1:0] matmul_16_och_count_buf;
  wire matmul_16_stream_pad_mask_0_0;
  assign matmul_16_stream_pad_mask_0_0 = (matmul_16_col_count + 0 < cparam_matmul_16_pad_col_left) || (matmul_16_col_count + 0 >= cparam_matmul_16_act_num_col + cparam_matmul_16_pad_col_left) || (matmul_16_row_count_buf + 0 < cparam_matmul_16_pad_row_top) || (matmul_16_row_count_buf + 0 >= cparam_matmul_16_act_num_row + cparam_matmul_16_pad_row_top);
  reg [1-1:0] matmul_16_stream_pad_masks;
  wire [14-1:0] stream_matmul_16_parameter_0_data;
  wire [1-1:0] stream_matmul_16_parameter_1_data;
  wire [1-1:0] stream_matmul_16_parameter_2_data;
  wire [1-1:0] stream_matmul_16_parameter_3_data;
  wire [2-1:0] stream_matmul_16_parameter_4_data;
  wire [1-1:0] stream_matmul_16__reduce_reset_data;
  wire [1-1:0] stream_matmul_16_parameter_6_data;
  wire [32-1:0] stream_matmul_16_source_7_data;
  wire [1-1:0] stream_matmul_16_parameter_8_data;
  wire [32-1:0] stream_matmul_16_source_9_data;
  wire [1-1:0] stream_matmul_16_parameter_10_data;
  wire [32-1:0] stream_matmul_16_source_11_data;
  wire [1-1:0] stream_matmul_16_parameter_12_data;
  wire [32-1:0] stream_matmul_16_source_13_data;
  wire [1-1:0] stream_matmul_16_parameter_14_data;
  wire [32-1:0] stream_matmul_16_source_15_data;
  wire [1-1:0] stream_matmul_16_parameter_16_data;
  wire [1-1:0] stream_matmul_16_parameter_17_data;
  wire [5-1:0] stream_matmul_16_parameter_18_data;
  wire [2-1:0] stream_matmul_16_parameter_19_data;
  wire [32-1:0] stream_matmul_16_source_20_data;
  wire [32-1:0] stream_matmul_16_source_21_data;
  wire [32-1:0] stream_matmul_16_source_22_data;
  reg __stream_matmul_16_stream_ivalid_1;
  reg __stream_matmul_16_stream_ivalid_2;
  reg __stream_matmul_16_stream_ivalid_3;
  reg __stream_matmul_16_stream_ivalid_4;
  reg __stream_matmul_16_stream_ivalid_5;
  reg __stream_matmul_16_stream_ivalid_6;
  reg __stream_matmul_16_stream_ivalid_7;
  reg __stream_matmul_16_stream_ivalid_8;
  reg __stream_matmul_16_stream_ivalid_9;
  reg __stream_matmul_16_stream_ivalid_10;
  reg __stream_matmul_16_stream_ivalid_11;
  reg __stream_matmul_16_stream_ivalid_12;
  reg __stream_matmul_16_stream_ivalid_13;
  reg __stream_matmul_16_stream_ivalid_14;
  reg __stream_matmul_16_stream_ivalid_15;
  reg __stream_matmul_16_stream_ivalid_16;
  reg __stream_matmul_16_stream_ivalid_17;
  reg __stream_matmul_16_stream_ivalid_18;
  reg __stream_matmul_16_stream_ivalid_19;
  reg __stream_matmul_16_stream_ivalid_20;
  reg __stream_matmul_16_stream_ivalid_21;
  reg __stream_matmul_16_stream_ivalid_22;
  reg __stream_matmul_16_stream_ivalid_23;
  reg __stream_matmul_16_stream_ivalid_24;
  reg __stream_matmul_16_stream_ivalid_25;
  reg __stream_matmul_16_stream_ivalid_26;
  reg __stream_matmul_16_stream_ivalid_27;
  reg __stream_matmul_16_stream_ivalid_28;
  reg __stream_matmul_16_stream_ivalid_29;
  reg __stream_matmul_16_stream_ivalid_30;
  reg __stream_matmul_16_stream_ivalid_31;
  reg __stream_matmul_16_stream_ivalid_32;
  reg [32-1:0] _counter_data_2451;
  reg [32-1:0] _counter_count_2451;
  wire _counter_reset_cond_2451;
  assign _counter_reset_cond_2451 = stream_matmul_16__reduce_reset_data;
  wire [32-1:0] _counter_current_count_2451;
  assign _counter_current_count_2451 = (_counter_reset_cond_2451)? 1'sd0 : _counter_count_2451;
  wire [1-1:0] _pointer_data_2454;
  assign _pointer_data_2454 = stream_matmul_16_parameter_4_data[1'sd0];
  reg [14-1:0] _minus_data_2456;
  wire [1-1:0] _pointer_data_2460;
  assign _pointer_data_2460 = stream_matmul_16_parameter_4_data[2'sd1];
  reg [14-1:0] _minus_data_2462;
  wire [16-1:0] _slice_data_2470;
  assign _slice_data_2470 = stream_matmul_16_source_7_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2471;
  assign _reinterpretcast_src_2471 = _slice_data_2470;
  wire signed [16-1:0] _reinterpretcast_data_2471;
  assign _reinterpretcast_data_2471 = _reinterpretcast_src_2471;
  wire [16-1:0] _slice_data_2474;
  assign _slice_data_2474 = stream_matmul_16_source_7_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2475;
  assign _reinterpretcast_src_2475 = _slice_data_2474;
  wire signed [16-1:0] _reinterpretcast_data_2475;
  assign _reinterpretcast_data_2475 = _reinterpretcast_src_2475;
  wire signed [16-1:0] _cond_data_2476;
  assign _cond_data_2476 = (stream_matmul_16_parameter_6_data)? _reinterpretcast_data_2471 : _reinterpretcast_data_2471;
  wire signed [16-1:0] _cond_data_2477;
  assign _cond_data_2477 = (stream_matmul_16_parameter_6_data)? _reinterpretcast_data_2471 : _reinterpretcast_data_2475;
  wire [16-1:0] _slice_data_2482;
  assign _slice_data_2482 = stream_matmul_16_source_9_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2483;
  assign _reinterpretcast_src_2483 = _slice_data_2482;
  wire signed [16-1:0] _reinterpretcast_data_2483;
  assign _reinterpretcast_data_2483 = _reinterpretcast_src_2483;
  wire [16-1:0] _slice_data_2486;
  assign _slice_data_2486 = stream_matmul_16_source_9_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2487;
  assign _reinterpretcast_src_2487 = _slice_data_2486;
  wire signed [16-1:0] _reinterpretcast_data_2487;
  assign _reinterpretcast_data_2487 = _reinterpretcast_src_2487;
  wire signed [16-1:0] _cond_data_2488;
  assign _cond_data_2488 = (stream_matmul_16_parameter_8_data)? _reinterpretcast_data_2483 : _reinterpretcast_data_2483;
  wire signed [16-1:0] _cond_data_2489;
  assign _cond_data_2489 = (stream_matmul_16_parameter_8_data)? _reinterpretcast_data_2483 : _reinterpretcast_data_2487;
  wire [16-1:0] _slice_data_2494;
  assign _slice_data_2494 = stream_matmul_16_source_11_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2495;
  assign _reinterpretcast_src_2495 = _slice_data_2494;
  wire [16-1:0] _reinterpretcast_data_2495;
  assign _reinterpretcast_data_2495 = _reinterpretcast_src_2495;
  wire [16-1:0] _slice_data_2498;
  assign _slice_data_2498 = stream_matmul_16_source_11_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2499;
  assign _reinterpretcast_src_2499 = _slice_data_2498;
  wire [16-1:0] _reinterpretcast_data_2499;
  assign _reinterpretcast_data_2499 = _reinterpretcast_src_2499;
  wire [16-1:0] _cond_data_2500;
  assign _cond_data_2500 = (stream_matmul_16_parameter_10_data)? _reinterpretcast_data_2495 : _reinterpretcast_data_2495;
  wire [16-1:0] _cond_data_2501;
  assign _cond_data_2501 = (stream_matmul_16_parameter_10_data)? _reinterpretcast_data_2495 : _reinterpretcast_data_2499;
  wire [16-1:0] _slice_data_2506;
  assign _slice_data_2506 = stream_matmul_16_source_13_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2507;
  assign _reinterpretcast_src_2507 = _slice_data_2506;
  wire [16-1:0] _reinterpretcast_data_2507;
  assign _reinterpretcast_data_2507 = _reinterpretcast_src_2507;
  wire [16-1:0] _slice_data_2510;
  assign _slice_data_2510 = stream_matmul_16_source_13_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2511;
  assign _reinterpretcast_src_2511 = _slice_data_2510;
  wire [16-1:0] _reinterpretcast_data_2511;
  assign _reinterpretcast_data_2511 = _reinterpretcast_src_2511;
  wire [16-1:0] _cond_data_2512;
  assign _cond_data_2512 = (stream_matmul_16_parameter_12_data)? _reinterpretcast_data_2507 : _reinterpretcast_data_2507;
  wire [16-1:0] _cond_data_2513;
  assign _cond_data_2513 = (stream_matmul_16_parameter_12_data)? _reinterpretcast_data_2507 : _reinterpretcast_data_2511;
  wire [16-1:0] _slice_data_2518;
  assign _slice_data_2518 = stream_matmul_16_source_15_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2519;
  assign _reinterpretcast_src_2519 = _slice_data_2518;
  wire [16-1:0] _reinterpretcast_data_2519;
  assign _reinterpretcast_data_2519 = _reinterpretcast_src_2519;
  wire [16-1:0] _slice_data_2522;
  assign _slice_data_2522 = stream_matmul_16_source_15_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2523;
  assign _reinterpretcast_src_2523 = _slice_data_2522;
  wire [16-1:0] _reinterpretcast_data_2523;
  assign _reinterpretcast_data_2523 = _reinterpretcast_src_2523;
  wire [16-1:0] _cond_data_2524;
  assign _cond_data_2524 = (stream_matmul_16_parameter_14_data)? _reinterpretcast_data_2519 : _reinterpretcast_data_2519;
  wire [16-1:0] _cond_data_2525;
  assign _cond_data_2525 = (stream_matmul_16_parameter_14_data)? _reinterpretcast_data_2519 : _reinterpretcast_data_2523;
  reg [1-1:0] _eq_data_2531;
  reg [1-1:0] _eq_data_2535;
  wire [16-1:0] _slice_data_2555;
  assign _slice_data_2555 = stream_matmul_16_source_21_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2556;
  assign _reinterpretcast_src_2556 = _slice_data_2555;
  wire signed [16-1:0] _reinterpretcast_data_2556;
  assign _reinterpretcast_data_2556 = _reinterpretcast_src_2556;
  wire [16-1:0] _slice_data_2559;
  assign _slice_data_2559 = stream_matmul_16_source_21_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2560;
  assign _reinterpretcast_src_2560 = _slice_data_2559;
  wire signed [16-1:0] _reinterpretcast_data_2560;
  assign _reinterpretcast_data_2560 = _reinterpretcast_src_2560;
  wire [16-1:0] _slice_data_2567;
  assign _slice_data_2567 = stream_matmul_16_source_22_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2568;
  assign _reinterpretcast_src_2568 = _slice_data_2567;
  wire signed [16-1:0] _reinterpretcast_data_2568;
  assign _reinterpretcast_data_2568 = _reinterpretcast_src_2568;
  wire [16-1:0] _slice_data_2571;
  assign _slice_data_2571 = stream_matmul_16_source_22_data[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2572;
  assign _reinterpretcast_src_2572 = _slice_data_2571;
  wire signed [16-1:0] _reinterpretcast_data_2572;
  assign _reinterpretcast_data_2572 = _reinterpretcast_src_2572;
  wire [1-1:0] _pointer_data_2577;
  assign _pointer_data_2577 = stream_matmul_16_parameter_3_data[1'sd0];
  reg [16-1:0] _plus_data_2582;
  reg [16-1:0] _plus_data_2587;
  reg [16-1:0] _plus_data_2592;
  reg [16-1:0] _plus_data_2597;
  reg [1-1:0] _eq_data_2603;
  reg [1-1:0] _eq_data_2606;
  reg [16-1:0] _plus_data_2613;
  reg [16-1:0] _plus_data_2618;
  reg [16-1:0] _plus_data_2623;
  reg [16-1:0] _plus_data_2628;
  reg [1-1:0] _eq_data_2634;
  reg [1-1:0] _eq_data_2637;
  reg [1-1:0] __delay_data_3119_pointer_2454;
  reg [32-1:0] __delay_data_3121__variable_2530;
  reg [1-1:0] __delay_data_3124_pointer_2577;
  reg signed [16-1:0] __delay_data_3127_reinterpretcast_2556;
  reg [1-1:0] __delay_data_3132_pointer_2460;
  reg signed [16-1:0] __delay_data_3136_reinterpretcast_2560;
  reg [1-1:0] __delay_data_3141__variable_2450;
  reg [14-1:0] __delay_data_3168__variable_2445;
  reg signed [16-1:0] __delay_data_3182_reinterpretcast_2568;
  reg signed [16-1:0] __delay_data_3187_reinterpretcast_2572;
  reg signed [16-1:0] __delay_data_3205_cond_2477;
  reg signed [16-1:0] __delay_data_3225_cond_2489;
  reg signed [16-1:0] __delay_data_3330_cond_2476;
  reg signed [16-1:0] __delay_data_3350_cond_2488;
  reg [1-1:0] _eq_data_2458;
  reg [1-1:0] _eq_data_2464;
  wire signed [32-1:0] _cond_data_2533;
  assign _cond_data_2533 = (_eq_data_2531)? __delay_data_3121__variable_2530 : 1'sd0;
  wire signed [32-1:0] _cond_data_2537;
  assign _cond_data_2537 = (_eq_data_2535)? _cond_data_2533 : 1'sd0;
  wire [16-1:0] _slice_data_2541;
  assign _slice_data_2541 = _cond_data_2537[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2542;
  assign _reinterpretcast_src_2542 = _slice_data_2541;
  wire signed [16-1:0] _reinterpretcast_data_2542;
  assign _reinterpretcast_data_2542 = _reinterpretcast_src_2542;
  wire [16-1:0] _slice_data_2545;
  assign _slice_data_2545 = _cond_data_2537[6'd31:6'd16];
  wire [16-1:0] _reinterpretcast_src_2546;
  assign _reinterpretcast_src_2546 = _slice_data_2545;
  wire signed [16-1:0] _reinterpretcast_data_2546;
  assign _reinterpretcast_data_2546 = _reinterpretcast_src_2546;
  reg [1-1:0] __delay_data_3120__delay_3119_pointer_2454;
  reg signed [16-1:0] __delay_data_3122_reinterpretcast_2542;
  reg [1-1:0] __delay_data_3125__delay_3124_pointer_2577;
  reg signed [16-1:0] __delay_data_3128__delay_3127_reinterpretcast_2556;
  reg [16-1:0] __delay_data_3130_plus_2582;
  reg [1-1:0] __delay_data_3133__delay_3132_pointer_2460;
  reg signed [16-1:0] __delay_data_3134_reinterpretcast_2546;
  reg signed [16-1:0] __delay_data_3137__delay_3136_reinterpretcast_2560;
  reg [16-1:0] __delay_data_3139_plus_2587;
  reg [1-1:0] __delay_data_3142__delay_3141__variable_2450;
  reg [16-1:0] __delay_data_3155_plus_2592;
  reg [14-1:0] __delay_data_3169__delay_3168__variable_2445;
  reg signed [16-1:0] __delay_data_3183__delay_3182_reinterpretcast_2568;
  reg [16-1:0] __delay_data_3185_plus_2613;
  reg signed [16-1:0] __delay_data_3188__delay_3187_reinterpretcast_2572;
  reg [16-1:0] __delay_data_3190_plus_2618;
  reg [16-1:0] __delay_data_3192_plus_2623;
  reg signed [16-1:0] __delay_data_3206__delay_3205_cond_2477;
  reg signed [16-1:0] __delay_data_3226__delay_3225_cond_2489;
  reg [16-1:0] __delay_data_3246_plus_2628;
  reg [1-1:0] __delay_data_3267_eq_2634;
  reg [1-1:0] __delay_data_3299_eq_2637;
  reg signed [16-1:0] __delay_data_3331__delay_3330_cond_2476;
  reg signed [16-1:0] __delay_data_3351__delay_3350_cond_2488;
  reg [16-1:0] __delay_data_3371_plus_2597;
  reg [1-1:0] __delay_data_3392_eq_2603;
  reg [1-1:0] __delay_data_3424_eq_2606;
  reg [1-1:0] _land_data_2459;
  reg [1-1:0] _land_data_2465;
  reg signed [16-1:0] __delay_data_3123__delay_3122_reinterpretcast_2542;
  reg [1-1:0] __delay_data_3126__delay_3125__delay_3124_pointer_2577;
  reg signed [16-1:0] __delay_data_3129__delay_3128__delay_3127_reinterpretcast_2556;
  reg [16-1:0] __delay_data_3131__delay_3130_plus_2582;
  reg signed [16-1:0] __delay_data_3135__delay_3134_reinterpretcast_2546;
  reg signed [16-1:0] __delay_data_3138__delay_3137__delay_3136_reinterpretcast_2560;
  reg [16-1:0] __delay_data_3140__delay_3139_plus_2587;
  reg [1-1:0] __delay_data_3143__delay_3142__delay_3141__variable_2450;
  reg [16-1:0] __delay_data_3156__delay_3155_plus_2592;
  reg [14-1:0] __delay_data_3170__delay_3169__delay_3168__variable_2445;
  reg signed [16-1:0] __delay_data_3184__delay_3183__delay_3182_reinterpretcast_2568;
  reg [16-1:0] __delay_data_3186__delay_3185_plus_2613;
  reg signed [16-1:0] __delay_data_3189__delay_3188__delay_3187_reinterpretcast_2572;
  reg [16-1:0] __delay_data_3191__delay_3190_plus_2618;
  reg [16-1:0] __delay_data_3193__delay_3192_plus_2623;
  reg signed [16-1:0] __delay_data_3207__delay_3206__delay_3205_cond_2477;
  reg signed [16-1:0] __delay_data_3227__delay_3226__delay_3225_cond_2489;
  reg [16-1:0] __delay_data_3247__delay_3246_plus_2628;
  reg [1-1:0] __delay_data_3268__delay_3267_eq_2634;
  reg [1-1:0] __delay_data_3300__delay_3299_eq_2637;
  reg signed [16-1:0] __delay_data_3332__delay_3331__delay_3330_cond_2476;
  reg signed [16-1:0] __delay_data_3352__delay_3351__delay_3350_cond_2488;
  reg [16-1:0] __delay_data_3372__delay_3371_plus_2597;
  reg [1-1:0] __delay_data_3393__delay_3392_eq_2603;
  reg [1-1:0] __delay_data_3425__delay_3424_eq_2606;
  wire signed [16-1:0] _cond_data_2548;
  assign _cond_data_2548 = (_land_data_2459)? 1'sd0 : __delay_data_3123__delay_3122_reinterpretcast_2542;
  wire signed [16-1:0] _cond_data_2550;
  assign _cond_data_2550 = (_land_data_2465)? 1'sd0 : __delay_data_3135__delay_3134_reinterpretcast_2546;
  wire signed [16-1:0] _cond_data_2562;
  assign _cond_data_2562 = (_land_data_2459)? 1'sd0 : __delay_data_3129__delay_3128__delay_3127_reinterpretcast_2556;
  wire signed [16-1:0] _cond_data_2564;
  assign _cond_data_2564 = (_land_data_2465)? 1'sd0 : __delay_data_3138__delay_3137__delay_3136_reinterpretcast_2560;
  wire signed [16-1:0] _cond_data_2574;
  assign _cond_data_2574 = (_land_data_2459)? 1'sd0 : __delay_data_3184__delay_3183__delay_3182_reinterpretcast_2568;
  wire signed [16-1:0] _cond_data_2576;
  assign _cond_data_2576 = (_land_data_2465)? 1'sd0 : __delay_data_3189__delay_3188__delay_3187_reinterpretcast_2572;
  wire signed [16-1:0] _cond_data_2580;
  assign _cond_data_2580 = (__delay_data_3126__delay_3125__delay_3124_pointer_2577)? 1'sd0 : _cond_data_2548;
  assign _mul_8_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_8_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_8_stream_internal_oready);
  wire signed [16-1:0] _cond_data_2585;
  assign _cond_data_2585 = (__delay_data_3126__delay_3125__delay_3124_pointer_2577)? 1'sd0 : _cond_data_2550;
  assign _mul_9_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_9_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_9_stream_internal_oready);
  wire signed [16-1:0] _cond_data_2611;
  assign _cond_data_2611 = (__delay_data_3126__delay_3125__delay_3124_pointer_2577)? 1'sd0 : _cond_data_2548;
  assign _mul_10_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_10_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_10_stream_internal_oready);
  wire signed [16-1:0] _cond_data_2616;
  assign _cond_data_2616 = (__delay_data_3126__delay_3125__delay_3124_pointer_2577)? 1'sd0 : _cond_data_2550;
  assign _mul_11_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_11_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_11_stream_internal_oready);
  reg [1-1:0] __delay_data_3144__delay_3143__delay_3142____variable_2450;
  reg [16-1:0] __delay_data_3157__delay_3156__delay_3155_plus_2592;
  reg [14-1:0] __delay_data_3171__delay_3170__delay_3169____variable_2445;
  reg [16-1:0] __delay_data_3194__delay_3193__delay_3192_plus_2623;
  reg signed [16-1:0] __delay_data_3208__delay_3207__delay_3206___cond_2477;
  reg signed [16-1:0] __delay_data_3228__delay_3227__delay_3226___cond_2489;
  reg [16-1:0] __delay_data_3248__delay_3247__delay_3246_plus_2628;
  reg [1-1:0] __delay_data_3269__delay_3268__delay_3267_eq_2634;
  reg [1-1:0] __delay_data_3301__delay_3300__delay_3299_eq_2637;
  reg signed [16-1:0] __delay_data_3333__delay_3332__delay_3331___cond_2476;
  reg signed [16-1:0] __delay_data_3353__delay_3352__delay_3351___cond_2488;
  reg [16-1:0] __delay_data_3373__delay_3372__delay_3371_plus_2597;
  reg [1-1:0] __delay_data_3394__delay_3393__delay_3392_eq_2603;
  reg [1-1:0] __delay_data_3426__delay_3425__delay_3424_eq_2606;
  reg [1-1:0] __delay_data_3145__delay_3144__delay_3143____variable_2450;
  reg [16-1:0] __delay_data_3158__delay_3157__delay_3156___plus_2592;
  reg [14-1:0] __delay_data_3172__delay_3171__delay_3170____variable_2445;
  reg [16-1:0] __delay_data_3195__delay_3194__delay_3193___plus_2623;
  reg signed [16-1:0] __delay_data_3209__delay_3208__delay_3207___cond_2477;
  reg signed [16-1:0] __delay_data_3229__delay_3228__delay_3227___cond_2489;
  reg [16-1:0] __delay_data_3249__delay_3248__delay_3247___plus_2628;
  reg [1-1:0] __delay_data_3270__delay_3269__delay_3268__delay_3267_eq_2634;
  reg [1-1:0] __delay_data_3302__delay_3301__delay_3300__delay_3299_eq_2637;
  reg signed [16-1:0] __delay_data_3334__delay_3333__delay_3332___cond_2476;
  reg signed [16-1:0] __delay_data_3354__delay_3353__delay_3352___cond_2488;
  reg [16-1:0] __delay_data_3374__delay_3373__delay_3372___plus_2597;
  reg [1-1:0] __delay_data_3395__delay_3394__delay_3393__delay_3392_eq_2603;
  reg [1-1:0] __delay_data_3427__delay_3426__delay_3425__delay_3424_eq_2606;
  reg [1-1:0] __delay_data_3146__delay_3145__delay_3144____variable_2450;
  reg [16-1:0] __delay_data_3159__delay_3158__delay_3157___plus_2592;
  reg [14-1:0] __delay_data_3173__delay_3172__delay_3171____variable_2445;
  reg [16-1:0] __delay_data_3196__delay_3195__delay_3194___plus_2623;
  reg signed [16-1:0] __delay_data_3210__delay_3209__delay_3208___cond_2477;
  reg signed [16-1:0] __delay_data_3230__delay_3229__delay_3228___cond_2489;
  reg [16-1:0] __delay_data_3250__delay_3249__delay_3248___plus_2628;
  reg [1-1:0] __delay_data_3271__delay_3270__delay_3269__delay_3268___eq_2634;
  reg [1-1:0] __delay_data_3303__delay_3302__delay_3301__delay_3300___eq_2637;
  reg signed [16-1:0] __delay_data_3335__delay_3334__delay_3333___cond_2476;
  reg signed [16-1:0] __delay_data_3355__delay_3354__delay_3353___cond_2488;
  reg [16-1:0] __delay_data_3375__delay_3374__delay_3373___plus_2597;
  reg [1-1:0] __delay_data_3396__delay_3395__delay_3394__delay_3393___eq_2603;
  reg [1-1:0] __delay_data_3428__delay_3427__delay_3426__delay_3425___eq_2606;
  reg [1-1:0] __delay_data_3147__delay_3146__delay_3145____variable_2450;
  reg [16-1:0] __delay_data_3160__delay_3159__delay_3158___plus_2592;
  reg [14-1:0] __delay_data_3174__delay_3173__delay_3172____variable_2445;
  reg [16-1:0] __delay_data_3197__delay_3196__delay_3195___plus_2623;
  reg signed [16-1:0] __delay_data_3211__delay_3210__delay_3209___cond_2477;
  reg signed [16-1:0] __delay_data_3231__delay_3230__delay_3229___cond_2489;
  reg [16-1:0] __delay_data_3251__delay_3250__delay_3249___plus_2628;
  reg [1-1:0] __delay_data_3272__delay_3271__delay_3270__delay_3269___eq_2634;
  reg [1-1:0] __delay_data_3304__delay_3303__delay_3302__delay_3301___eq_2637;
  reg signed [16-1:0] __delay_data_3336__delay_3335__delay_3334___cond_2476;
  reg signed [16-1:0] __delay_data_3356__delay_3355__delay_3354___cond_2488;
  reg [16-1:0] __delay_data_3376__delay_3375__delay_3374___plus_2597;
  reg [1-1:0] __delay_data_3397__delay_3396__delay_3395__delay_3394___eq_2603;
  reg [1-1:0] __delay_data_3429__delay_3428__delay_3427__delay_3426___eq_2606;
  reg [1-1:0] __delay_data_3148__delay_3147__delay_3146____variable_2450;
  reg [16-1:0] __delay_data_3161__delay_3160__delay_3159___plus_2592;
  reg [14-1:0] __delay_data_3175__delay_3174__delay_3173____variable_2445;
  reg [16-1:0] __delay_data_3198__delay_3197__delay_3196___plus_2623;
  reg signed [16-1:0] __delay_data_3212__delay_3211__delay_3210___cond_2477;
  reg signed [16-1:0] __delay_data_3232__delay_3231__delay_3230___cond_2489;
  reg [16-1:0] __delay_data_3252__delay_3251__delay_3250___plus_2628;
  reg [1-1:0] __delay_data_3273__delay_3272__delay_3271__delay_3270___eq_2634;
  reg [1-1:0] __delay_data_3305__delay_3304__delay_3303__delay_3302___eq_2637;
  reg signed [16-1:0] __delay_data_3337__delay_3336__delay_3335___cond_2476;
  reg signed [16-1:0] __delay_data_3357__delay_3356__delay_3355___cond_2488;
  reg [16-1:0] __delay_data_3377__delay_3376__delay_3375___plus_2597;
  reg [1-1:0] __delay_data_3398__delay_3397__delay_3396__delay_3395___eq_2603;
  reg [1-1:0] __delay_data_3430__delay_3429__delay_3428__delay_3427___eq_2606;
  reg [1-1:0] __delay_data_3149__delay_3148__delay_3147____variable_2450;
  reg [16-1:0] __delay_data_3162__delay_3161__delay_3160___plus_2592;
  reg [14-1:0] __delay_data_3176__delay_3175__delay_3174____variable_2445;
  reg [16-1:0] __delay_data_3199__delay_3198__delay_3197___plus_2623;
  reg signed [16-1:0] __delay_data_3213__delay_3212__delay_3211___cond_2477;
  reg signed [16-1:0] __delay_data_3233__delay_3232__delay_3231___cond_2489;
  reg [16-1:0] __delay_data_3253__delay_3252__delay_3251___plus_2628;
  reg [1-1:0] __delay_data_3274__delay_3273__delay_3272__delay_3271___eq_2634;
  reg [1-1:0] __delay_data_3306__delay_3305__delay_3304__delay_3303___eq_2637;
  reg signed [16-1:0] __delay_data_3338__delay_3337__delay_3336___cond_2476;
  reg signed [16-1:0] __delay_data_3358__delay_3357__delay_3356___cond_2488;
  reg [16-1:0] __delay_data_3378__delay_3377__delay_3376___plus_2597;
  reg [1-1:0] __delay_data_3399__delay_3398__delay_3397__delay_3396___eq_2603;
  reg [1-1:0] __delay_data_3431__delay_3430__delay_3429__delay_3428___eq_2606;
  reg [1-1:0] __delay_data_3150__delay_3149__delay_3148____variable_2450;
  reg [16-1:0] __delay_data_3163__delay_3162__delay_3161___plus_2592;
  reg [14-1:0] __delay_data_3177__delay_3176__delay_3175____variable_2445;
  reg [16-1:0] __delay_data_3200__delay_3199__delay_3198___plus_2623;
  reg signed [16-1:0] __delay_data_3214__delay_3213__delay_3212___cond_2477;
  reg signed [16-1:0] __delay_data_3234__delay_3233__delay_3232___cond_2489;
  reg [16-1:0] __delay_data_3254__delay_3253__delay_3252___plus_2628;
  reg [1-1:0] __delay_data_3275__delay_3274__delay_3273__delay_3272___eq_2634;
  reg [1-1:0] __delay_data_3307__delay_3306__delay_3305__delay_3304___eq_2637;
  reg signed [16-1:0] __delay_data_3339__delay_3338__delay_3337___cond_2476;
  reg signed [16-1:0] __delay_data_3359__delay_3358__delay_3357___cond_2488;
  reg [16-1:0] __delay_data_3379__delay_3378__delay_3377___plus_2597;
  reg [1-1:0] __delay_data_3400__delay_3399__delay_3398__delay_3397___eq_2603;
  reg [1-1:0] __delay_data_3432__delay_3431__delay_3430__delay_3429___eq_2606;
  reg [1-1:0] __delay_data_3151__delay_3150__delay_3149____variable_2450;
  reg [16-1:0] __delay_data_3164__delay_3163__delay_3162___plus_2592;
  reg [14-1:0] __delay_data_3178__delay_3177__delay_3176____variable_2445;
  reg [16-1:0] __delay_data_3201__delay_3200__delay_3199___plus_2623;
  reg signed [16-1:0] __delay_data_3215__delay_3214__delay_3213___cond_2477;
  reg signed [16-1:0] __delay_data_3235__delay_3234__delay_3233___cond_2489;
  reg [16-1:0] __delay_data_3255__delay_3254__delay_3253___plus_2628;
  reg [1-1:0] __delay_data_3276__delay_3275__delay_3274__delay_3273___eq_2634;
  reg [1-1:0] __delay_data_3308__delay_3307__delay_3306__delay_3305___eq_2637;
  reg signed [16-1:0] __delay_data_3340__delay_3339__delay_3338___cond_2476;
  reg signed [16-1:0] __delay_data_3360__delay_3359__delay_3358___cond_2488;
  reg [16-1:0] __delay_data_3380__delay_3379__delay_3378___plus_2597;
  reg [1-1:0] __delay_data_3401__delay_3400__delay_3399__delay_3398___eq_2603;
  reg [1-1:0] __delay_data_3433__delay_3432__delay_3431__delay_3430___eq_2606;
  reg [1-1:0] __delay_data_3152__delay_3151__delay_3150____variable_2450;
  reg [16-1:0] __delay_data_3165__delay_3164__delay_3163___plus_2592;
  reg [14-1:0] __delay_data_3179__delay_3178__delay_3177____variable_2445;
  reg [16-1:0] __delay_data_3202__delay_3201__delay_3200___plus_2623;
  reg signed [16-1:0] __delay_data_3216__delay_3215__delay_3214___cond_2477;
  reg signed [16-1:0] __delay_data_3236__delay_3235__delay_3234___cond_2489;
  reg [16-1:0] __delay_data_3256__delay_3255__delay_3254___plus_2628;
  reg [1-1:0] __delay_data_3277__delay_3276__delay_3275__delay_3274___eq_2634;
  reg [1-1:0] __delay_data_3309__delay_3308__delay_3307__delay_3306___eq_2637;
  reg signed [16-1:0] __delay_data_3341__delay_3340__delay_3339___cond_2476;
  reg signed [16-1:0] __delay_data_3361__delay_3360__delay_3359___cond_2488;
  reg [16-1:0] __delay_data_3381__delay_3380__delay_3379___plus_2597;
  reg [1-1:0] __delay_data_3402__delay_3401__delay_3400__delay_3399___eq_2603;
  reg [1-1:0] __delay_data_3434__delay_3433__delay_3432__delay_3431___eq_2606;
  wire signed [32-1:0] __substreamoutput_data_2583;
  assign __substreamoutput_data_2583 = mul_8_z_data;
  wire signed [32-1:0] __substreamoutput_data_2588;
  assign __substreamoutput_data_2588 = mul_9_z_data;
  reg signed [64-1:0] __variable_wdata_44;
  assign add_tree_2_var0_data = __variable_wdata_44;
  reg signed [64-1:0] __variable_wdata_45;
  assign add_tree_2_var1_data = __variable_wdata_45;
  assign _add_tree_2_is_root = ((_stream_matmul_16_busy)? 0 : 1) && 1;
  assign _add_tree_2_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && _add_tree_2_stream_internal_oready;
  wire signed [32-1:0] __substreamoutput_data_2614;
  assign __substreamoutput_data_2614 = mul_10_z_data;
  wire signed [32-1:0] __substreamoutput_data_2619;
  assign __substreamoutput_data_2619 = mul_11_z_data;
  reg signed [64-1:0] __variable_wdata_48;
  assign add_tree_3_var0_data = __variable_wdata_48;
  reg signed [64-1:0] __variable_wdata_49;
  assign add_tree_3_var1_data = __variable_wdata_49;
  assign _add_tree_3_is_root = ((_stream_matmul_16_busy)? 0 : 1) && 1;
  assign _add_tree_3_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && _add_tree_3_stream_internal_oready;
  reg [1-1:0] __delay_data_3153__delay_3152__delay_3151____variable_2450;
  reg [16-1:0] __delay_data_3166__delay_3165__delay_3164___plus_2592;
  reg [14-1:0] __delay_data_3180__delay_3179__delay_3178____variable_2445;
  reg [16-1:0] __delay_data_3203__delay_3202__delay_3201___plus_2623;
  reg signed [16-1:0] __delay_data_3217__delay_3216__delay_3215___cond_2477;
  reg signed [16-1:0] __delay_data_3237__delay_3236__delay_3235___cond_2489;
  reg [16-1:0] __delay_data_3257__delay_3256__delay_3255___plus_2628;
  reg [1-1:0] __delay_data_3278__delay_3277__delay_3276__delay_3275___eq_2634;
  reg [1-1:0] __delay_data_3310__delay_3309__delay_3308__delay_3307___eq_2637;
  reg signed [16-1:0] __delay_data_3342__delay_3341__delay_3340___cond_2476;
  reg signed [16-1:0] __delay_data_3362__delay_3361__delay_3360___cond_2488;
  reg [16-1:0] __delay_data_3382__delay_3381__delay_3380___plus_2597;
  reg [1-1:0] __delay_data_3403__delay_3402__delay_3401__delay_3400___eq_2603;
  reg [1-1:0] __delay_data_3435__delay_3434__delay_3433__delay_3432___eq_2606;
  reg [1-1:0] __delay_data_3154__delay_3153__delay_3152____variable_2450;
  reg [16-1:0] __delay_data_3167__delay_3166__delay_3165___plus_2592;
  reg [14-1:0] __delay_data_3181__delay_3180__delay_3179____variable_2445;
  reg [16-1:0] __delay_data_3204__delay_3203__delay_3202___plus_2623;
  reg signed [16-1:0] __delay_data_3218__delay_3217__delay_3216___cond_2477;
  reg signed [16-1:0] __delay_data_3238__delay_3237__delay_3236___cond_2489;
  reg [16-1:0] __delay_data_3258__delay_3257__delay_3256___plus_2628;
  reg [1-1:0] __delay_data_3279__delay_3278__delay_3277__delay_3276___eq_2634;
  reg [1-1:0] __delay_data_3311__delay_3310__delay_3309__delay_3308___eq_2637;
  reg signed [16-1:0] __delay_data_3343__delay_3342__delay_3341___cond_2476;
  reg signed [16-1:0] __delay_data_3363__delay_3362__delay_3361___cond_2488;
  reg [16-1:0] __delay_data_3383__delay_3382__delay_3381___plus_2597;
  reg [1-1:0] __delay_data_3404__delay_3403__delay_3402__delay_3401___eq_2603;
  reg [1-1:0] __delay_data_3436__delay_3435__delay_3434__delay_3433___eq_2606;
  wire signed [64-1:0] __substreamoutput_data_2590;
  assign __substreamoutput_data_2590 = add_tree_2_sum_data;
  assign _acc_0_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _acc_0_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _acc_0_stream_internal_oready);
  wire signed [64-1:0] __substreamoutput_data_2621;
  assign __substreamoutput_data_2621 = add_tree_3_sum_data;
  assign _acc_1_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _acc_1_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _acc_1_stream_internal_oready);
  reg signed [16-1:0] __delay_data_3219__delay_3218__delay_3217___cond_2477;
  reg signed [16-1:0] __delay_data_3239__delay_3238__delay_3237___cond_2489;
  reg [16-1:0] __delay_data_3259__delay_3258__delay_3257___plus_2628;
  reg [1-1:0] __delay_data_3280__delay_3279__delay_3278__delay_3277___eq_2634;
  reg [1-1:0] __delay_data_3312__delay_3311__delay_3310__delay_3309___eq_2637;
  reg signed [16-1:0] __delay_data_3344__delay_3343__delay_3342___cond_2476;
  reg signed [16-1:0] __delay_data_3364__delay_3363__delay_3362___cond_2488;
  reg [16-1:0] __delay_data_3384__delay_3383__delay_3382___plus_2597;
  reg [1-1:0] __delay_data_3405__delay_3404__delay_3403__delay_3402___eq_2603;
  reg [1-1:0] __delay_data_3437__delay_3436__delay_3435__delay_3434___eq_2606;
  reg signed [16-1:0] __delay_data_3220__delay_3219__delay_3218___cond_2477;
  reg signed [16-1:0] __delay_data_3240__delay_3239__delay_3238___cond_2489;
  reg [16-1:0] __delay_data_3260__delay_3259__delay_3258___plus_2628;
  reg [1-1:0] __delay_data_3281__delay_3280__delay_3279__delay_3278___eq_2634;
  reg [1-1:0] __delay_data_3313__delay_3312__delay_3311__delay_3310___eq_2637;
  reg signed [16-1:0] __delay_data_3345__delay_3344__delay_3343___cond_2476;
  reg signed [16-1:0] __delay_data_3365__delay_3364__delay_3363___cond_2488;
  reg [16-1:0] __delay_data_3385__delay_3384__delay_3383___plus_2597;
  reg [1-1:0] __delay_data_3406__delay_3405__delay_3404__delay_3403___eq_2603;
  reg [1-1:0] __delay_data_3438__delay_3437__delay_3436__delay_3435___eq_2606;
  reg signed [16-1:0] __delay_data_3221__delay_3220__delay_3219___cond_2477;
  reg signed [16-1:0] __delay_data_3241__delay_3240__delay_3239___cond_2489;
  reg [16-1:0] __delay_data_3261__delay_3260__delay_3259___plus_2628;
  reg [1-1:0] __delay_data_3282__delay_3281__delay_3280__delay_3279___eq_2634;
  reg [1-1:0] __delay_data_3314__delay_3313__delay_3312__delay_3311___eq_2637;
  reg signed [16-1:0] __delay_data_3346__delay_3345__delay_3344___cond_2476;
  reg signed [16-1:0] __delay_data_3366__delay_3365__delay_3364___cond_2488;
  reg [16-1:0] __delay_data_3386__delay_3385__delay_3384___plus_2597;
  reg [1-1:0] __delay_data_3407__delay_3406__delay_3405__delay_3404___eq_2603;
  reg [1-1:0] __delay_data_3439__delay_3438__delay_3437__delay_3436___eq_2606;
  reg signed [16-1:0] __delay_data_3222__delay_3221__delay_3220___cond_2477;
  reg signed [16-1:0] __delay_data_3242__delay_3241__delay_3240___cond_2489;
  reg [16-1:0] __delay_data_3262__delay_3261__delay_3260___plus_2628;
  reg [1-1:0] __delay_data_3283__delay_3282__delay_3281__delay_3280___eq_2634;
  reg [1-1:0] __delay_data_3315__delay_3314__delay_3313__delay_3312___eq_2637;
  reg signed [16-1:0] __delay_data_3347__delay_3346__delay_3345___cond_2476;
  reg signed [16-1:0] __delay_data_3367__delay_3366__delay_3365___cond_2488;
  reg [16-1:0] __delay_data_3387__delay_3386__delay_3385___plus_2597;
  reg [1-1:0] __delay_data_3408__delay_3407__delay_3406__delay_3405___eq_2603;
  reg [1-1:0] __delay_data_3440__delay_3439__delay_3438__delay_3437___eq_2606;
  reg signed [16-1:0] __delay_data_3223__delay_3222__delay_3221___cond_2477;
  reg signed [16-1:0] __delay_data_3243__delay_3242__delay_3241___cond_2489;
  reg [16-1:0] __delay_data_3263__delay_3262__delay_3261___plus_2628;
  reg [1-1:0] __delay_data_3284__delay_3283__delay_3282__delay_3281___eq_2634;
  reg [1-1:0] __delay_data_3316__delay_3315__delay_3314__delay_3313___eq_2637;
  reg signed [16-1:0] __delay_data_3348__delay_3347__delay_3346___cond_2476;
  reg signed [16-1:0] __delay_data_3368__delay_3367__delay_3366___cond_2488;
  reg [16-1:0] __delay_data_3388__delay_3387__delay_3386___plus_2597;
  reg [1-1:0] __delay_data_3409__delay_3408__delay_3407__delay_3406___eq_2603;
  reg [1-1:0] __delay_data_3441__delay_3440__delay_3439__delay_3438___eq_2606;
  reg signed [16-1:0] __delay_data_3224__delay_3223__delay_3222___cond_2477;
  reg signed [16-1:0] __delay_data_3244__delay_3243__delay_3242___cond_2489;
  reg [16-1:0] __delay_data_3264__delay_3263__delay_3262___plus_2628;
  reg [1-1:0] __delay_data_3285__delay_3284__delay_3283__delay_3282___eq_2634;
  reg [1-1:0] __delay_data_3317__delay_3316__delay_3315__delay_3314___eq_2637;
  reg signed [16-1:0] __delay_data_3349__delay_3348__delay_3347___cond_2476;
  reg signed [16-1:0] __delay_data_3369__delay_3368__delay_3367___cond_2488;
  reg [16-1:0] __delay_data_3389__delay_3388__delay_3387___plus_2597;
  reg [1-1:0] __delay_data_3410__delay_3409__delay_3408__delay_3407___eq_2603;
  reg [1-1:0] __delay_data_3442__delay_3441__delay_3440__delay_3439___eq_2606;
  wire signed [64-1:0] __substreamoutput_data_2593;
  assign __substreamoutput_data_2593 = acc_0_sum_data;
  wire [1-1:0] __substreamoutput_data_2594;
  assign __substreamoutput_data_2594 = acc_0_valid_data;
  reg signed [64-1:0] _plus_data_2595;
  wire signed [64-1:0] __substreamoutput_data_2624;
  assign __substreamoutput_data_2624 = acc_1_sum_data;
  reg signed [64-1:0] _plus_data_2626;
  reg signed [16-1:0] __delay_data_3245__delay_3244__delay_3243___cond_2489;
  reg [16-1:0] __delay_data_3265__delay_3264__delay_3263___plus_2628;
  reg [1-1:0] __delay_data_3286__delay_3285__delay_3284__delay_3283___eq_2634;
  reg [1-1:0] __delay_data_3318__delay_3317__delay_3316__delay_3315___eq_2637;
  reg signed [16-1:0] __delay_data_3370__delay_3369__delay_3368___cond_2488;
  reg [16-1:0] __delay_data_3390__delay_3389__delay_3388___plus_2597;
  reg [1-1:0] __delay_data_3411__delay_3410__delay_3409__delay_3408___eq_2603;
  reg [1-1:0] __delay_data_3443__delay_3442__delay_3441__delay_3440___eq_2606;
  reg [1-1:0] __delay_data_3455__substreamoutput_2594;
  assign _mul_rshift_round_clip_6_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_rshift_round_clip_6_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_rshift_round_clip_6_stream_internal_oready);
  assign _mul_rshift_round_clip_7_is_root = ((_stream_matmul_16_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_rshift_round_clip_7_stream_oready = ((_stream_matmul_16_busy)? _stream_matmul_16_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_rshift_round_clip_7_stream_internal_oready);
  assign _stream_matmul_16_stream_internal_oready = ((_stream_matmul_16_busy)? _mul_rshift_round_clip_7_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _mul_rshift_round_clip_6_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _acc_1_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _acc_0_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _add_tree_3_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _add_tree_2_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _mul_11_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _mul_10_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _mul_9_stream_internal_oready : 1) && (((_stream_matmul_16_busy)? _mul_8_stream_internal_oready : 1) && 1)))))))));
  reg [1-1:0] __delay_data_3287__delay_3286__delay_3285__delay_3284___eq_2634;
  reg [1-1:0] __delay_data_3319__delay_3318__delay_3317__delay_3316___eq_2637;
  reg [1-1:0] __delay_data_3412__delay_3411__delay_3410__delay_3409___eq_2603;
  reg [1-1:0] __delay_data_3444__delay_3443__delay_3442__delay_3441___eq_2606;
  reg [1-1:0] __delay_data_3456__delay_3455__substreamoutput_2594;
  reg [1-1:0] __delay_data_3288__delay_3287__delay_3286__delay_3285___eq_2634;
  reg [1-1:0] __delay_data_3320__delay_3319__delay_3318__delay_3317___eq_2637;
  reg [1-1:0] __delay_data_3413__delay_3412__delay_3411__delay_3410___eq_2603;
  reg [1-1:0] __delay_data_3445__delay_3444__delay_3443__delay_3442___eq_2606;
  reg [1-1:0] __delay_data_3457__delay_3456____substreamoutput_2594;
  reg [1-1:0] __delay_data_3289__delay_3288__delay_3287__delay_3286___eq_2634;
  reg [1-1:0] __delay_data_3321__delay_3320__delay_3319__delay_3318___eq_2637;
  reg [1-1:0] __delay_data_3414__delay_3413__delay_3412__delay_3411___eq_2603;
  reg [1-1:0] __delay_data_3446__delay_3445__delay_3444__delay_3443___eq_2606;
  reg [1-1:0] __delay_data_3458__delay_3457____substreamoutput_2594;
  reg [1-1:0] __delay_data_3290__delay_3289__delay_3288__delay_3287___eq_2634;
  reg [1-1:0] __delay_data_3322__delay_3321__delay_3320__delay_3319___eq_2637;
  reg [1-1:0] __delay_data_3415__delay_3414__delay_3413__delay_3412___eq_2603;
  reg [1-1:0] __delay_data_3447__delay_3446__delay_3445__delay_3444___eq_2606;
  reg [1-1:0] __delay_data_3459__delay_3458____substreamoutput_2594;
  reg [1-1:0] __delay_data_3291__delay_3290__delay_3289__delay_3288___eq_2634;
  reg [1-1:0] __delay_data_3323__delay_3322__delay_3321__delay_3320___eq_2637;
  reg [1-1:0] __delay_data_3416__delay_3415__delay_3414__delay_3413___eq_2603;
  reg [1-1:0] __delay_data_3448__delay_3447__delay_3446__delay_3445___eq_2606;
  reg [1-1:0] __delay_data_3460__delay_3459____substreamoutput_2594;
  reg [1-1:0] __delay_data_3292__delay_3291__delay_3290__delay_3289___eq_2634;
  reg [1-1:0] __delay_data_3324__delay_3323__delay_3322__delay_3321___eq_2637;
  reg [1-1:0] __delay_data_3417__delay_3416__delay_3415__delay_3414___eq_2603;
  reg [1-1:0] __delay_data_3449__delay_3448__delay_3447__delay_3446___eq_2606;
  reg [1-1:0] __delay_data_3461__delay_3460____substreamoutput_2594;
  reg [1-1:0] __delay_data_3293__delay_3292__delay_3291__delay_3290___eq_2634;
  reg [1-1:0] __delay_data_3325__delay_3324__delay_3323__delay_3322___eq_2637;
  reg [1-1:0] __delay_data_3418__delay_3417__delay_3416__delay_3415___eq_2603;
  reg [1-1:0] __delay_data_3450__delay_3449__delay_3448__delay_3447___eq_2606;
  reg [1-1:0] __delay_data_3462__delay_3461____substreamoutput_2594;
  reg [1-1:0] __delay_data_3294__delay_3293__delay_3292__delay_3291___eq_2634;
  reg [1-1:0] __delay_data_3326__delay_3325__delay_3324__delay_3323___eq_2637;
  reg [1-1:0] __delay_data_3419__delay_3418__delay_3417__delay_3416___eq_2603;
  reg [1-1:0] __delay_data_3451__delay_3450__delay_3449__delay_3448___eq_2606;
  reg [1-1:0] __delay_data_3463__delay_3462____substreamoutput_2594;
  reg [1-1:0] __delay_data_3295__delay_3294__delay_3293__delay_3292___eq_2634;
  reg [1-1:0] __delay_data_3327__delay_3326__delay_3325__delay_3324___eq_2637;
  reg [1-1:0] __delay_data_3420__delay_3419__delay_3418__delay_3417___eq_2603;
  reg [1-1:0] __delay_data_3452__delay_3451__delay_3450__delay_3449___eq_2606;
  reg [1-1:0] __delay_data_3464__delay_3463____substreamoutput_2594;
  wire signed [16-1:0] __substreamoutput_data_2598;
  assign __substreamoutput_data_2598 = mul_rshift_round_clip_6_z_data;
  reg [1-1:0] _greaterthan_data_2600;
  wire signed [16-1:0] __substreamoutput_data_2629;
  assign __substreamoutput_data_2629 = mul_rshift_round_clip_7_z_data;
  reg [1-1:0] _greaterthan_data_2631;
  reg signed [16-1:0] __delay_data_3266__substreamoutput_2629;
  reg [1-1:0] __delay_data_3296__delay_3295__delay_3294__delay_3293___eq_2634;
  reg [1-1:0] __delay_data_3328__delay_3327__delay_3326__delay_3325___eq_2637;
  reg signed [16-1:0] __delay_data_3391__substreamoutput_2598;
  reg [1-1:0] __delay_data_3421__delay_3420__delay_3419__delay_3418___eq_2603;
  reg [1-1:0] __delay_data_3453__delay_3452__delay_3451__delay_3450___eq_2606;
  reg [1-1:0] __delay_data_3465__delay_3464____substreamoutput_2594;
  reg signed [16-1:0] _cond_data_2602;
  reg signed [16-1:0] _cond_data_2633;
  reg [1-1:0] __delay_data_3297__delay_3296__delay_3295__delay_3294___eq_2634;
  reg signed [16-1:0] __delay_data_3298__delay_3266__substreamoutput_2629;
  reg [1-1:0] __delay_data_3329__delay_3328__delay_3327__delay_3326___eq_2637;
  reg [1-1:0] __delay_data_3422__delay_3421__delay_3420__delay_3419___eq_2603;
  reg signed [16-1:0] __delay_data_3423__delay_3391__substreamoutput_2598;
  reg [1-1:0] __delay_data_3454__delay_3453__delay_3452__delay_3451___eq_2606;
  reg [1-1:0] __delay_data_3466__delay_3465____substreamoutput_2594;
  wire signed [16-1:0] _cond_data_2605;
  assign _cond_data_2605 = (__delay_data_3422__delay_3421__delay_3420__delay_3419___eq_2603)? _cond_data_2602 : __delay_data_3423__delay_3391__substreamoutput_2598;
  wire signed [16-1:0] _cond_data_2608;
  assign _cond_data_2608 = (__delay_data_3454__delay_3453__delay_3452__delay_3451___eq_2606)? __delay_data_3423__delay_3391__substreamoutput_2598 : _cond_data_2605;
  wire signed [16-1:0] _reinterpretcast_src_2609;
  assign _reinterpretcast_src_2609 = _cond_data_2608;
  wire signed [16-1:0] _reinterpretcast_data_2609;
  assign _reinterpretcast_data_2609 = _reinterpretcast_src_2609;
  wire signed [16-1:0] _cond_data_2636;
  assign _cond_data_2636 = (__delay_data_3297__delay_3296__delay_3295__delay_3294___eq_2634)? _cond_data_2633 : __delay_data_3298__delay_3266__substreamoutput_2629;
  wire signed [16-1:0] _cond_data_2639;
  assign _cond_data_2639 = (__delay_data_3329__delay_3328__delay_3327__delay_3326___eq_2637)? __delay_data_3298__delay_3266__substreamoutput_2629 : _cond_data_2636;
  wire signed [16-1:0] _reinterpretcast_src_2640;
  assign _reinterpretcast_src_2640 = _cond_data_2639;
  wire signed [16-1:0] _reinterpretcast_data_2640;
  assign _reinterpretcast_data_2640 = _reinterpretcast_src_2640;
  wire [32-1:0] _cat_data_2641;
  assign _cat_data_2641 = { _reinterpretcast_data_2640, _reinterpretcast_data_2609 };
  wire [32-1:0] stream_matmul_16_sink_33_data;
  assign stream_matmul_16_sink_33_data = _cat_data_2641;
  wire [1-1:0] stream_matmul_16_sink_34_data;
  assign stream_matmul_16_sink_34_data = __delay_data_3466__delay_3465____substreamoutput_2594;
  wire _set_flag_2207;
  assign _set_flag_2207 = matmul_16_comp_fsm == 3;
  reg [14-1:0] __variable_wdata_2445;
  assign stream_matmul_16_parameter_0_data = __variable_wdata_2445;
  wire _set_flag_2208;
  assign _set_flag_2208 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2446;
  assign stream_matmul_16_parameter_1_data = __variable_wdata_2446;
  wire _set_flag_2209;
  assign _set_flag_2209 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2447;
  assign stream_matmul_16_parameter_2_data = __variable_wdata_2447;
  wire _set_flag_2210;
  assign _set_flag_2210 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2448;
  assign stream_matmul_16_parameter_3_data = __variable_wdata_2448;
  wire _set_flag_2211;
  assign _set_flag_2211 = matmul_16_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_2449;
  assign stream_matmul_16_parameter_4_data = __variable_wdata_2449;
  wire _set_flag_2212;
  assign _set_flag_2212 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2466;
  assign stream_matmul_16_parameter_6_data = __variable_wdata_2466;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_0;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_1;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_2;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_3;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_count_0;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_count_1;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_count_2;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_count_3;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_16_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_16_source_7_pat_stride_buf_3;
  wire _set_flag_2213;
  assign _set_flag_2213 = matmul_16_comp_fsm == 3;
  assign ram_w32_l256_id0_0_addr = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_7_source_ram_renable && (_stream_matmul_16_source_7_source_sel == 1))? _stream_matmul_16_source_7_source_ram_raddr : 'hx;
  assign ram_w32_l256_id0_0_enable = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_7_source_ram_renable && (_stream_matmul_16_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_2214 = 1;
  wire [_tmp_2214-1:0] _tmp_2215;
  assign _tmp_2215 = _stream_matmul_16_stream_oready && _stream_matmul_16_source_7_source_ram_renable && (_stream_matmul_16_source_7_source_sel == 1);
  reg [_tmp_2214-1:0] __tmp_2215_1;
  assign _stream_matmul_16_source_7_source_ram_rdata = (_stream_matmul_16_source_7_source_sel == 1)? ram_w32_l256_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_2467;
  assign stream_matmul_16_source_7_data = __variable_wdata_2467;
  reg [32-1:0] _stream_matmul_16_source_7_source_pat_fsm_0;
  localparam _stream_matmul_16_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_matmul_16_source_7_source_pat_all_offset;
  assign _stream_matmul_16_source_7_source_pat_all_offset = _stream_matmul_16_source_7_source_offset_buf + _source_stream_matmul_16_source_7_pat_cur_offset_0 + _source_stream_matmul_16_source_7_pat_cur_offset_1 + _source_stream_matmul_16_source_7_pat_cur_offset_2 + _source_stream_matmul_16_source_7_pat_cur_offset_3;
  wire _set_flag_2216;
  assign _set_flag_2216 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2478;
  assign stream_matmul_16_parameter_8_data = __variable_wdata_2478;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_0;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_1;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_2;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_3;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_count_0;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_count_1;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_count_2;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_count_3;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_16_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_16_source_9_pat_stride_buf_3;
  wire _set_flag_2217;
  assign _set_flag_2217 = matmul_16_comp_fsm == 3;
  assign ram_w32_l256_id1_0_addr = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_9_source_ram_renable && (_stream_matmul_16_source_9_source_sel == 2))? _stream_matmul_16_source_9_source_ram_raddr : 'hx;
  assign ram_w32_l256_id1_0_enable = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_9_source_ram_renable && (_stream_matmul_16_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_2218 = 1;
  wire [_tmp_2218-1:0] _tmp_2219;
  assign _tmp_2219 = _stream_matmul_16_stream_oready && _stream_matmul_16_source_9_source_ram_renable && (_stream_matmul_16_source_9_source_sel == 2);
  reg [_tmp_2218-1:0] __tmp_2219_1;
  assign _stream_matmul_16_source_9_source_ram_rdata = (_stream_matmul_16_source_9_source_sel == 2)? ram_w32_l256_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_2479;
  assign stream_matmul_16_source_9_data = __variable_wdata_2479;
  reg [32-1:0] _stream_matmul_16_source_9_source_pat_fsm_1;
  localparam _stream_matmul_16_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_matmul_16_source_9_source_pat_all_offset;
  assign _stream_matmul_16_source_9_source_pat_all_offset = _stream_matmul_16_source_9_source_offset_buf + _source_stream_matmul_16_source_9_pat_cur_offset_0 + _source_stream_matmul_16_source_9_pat_cur_offset_1 + _source_stream_matmul_16_source_9_pat_cur_offset_2 + _source_stream_matmul_16_source_9_pat_cur_offset_3;
  wire _set_flag_2220;
  assign _set_flag_2220 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2490;
  assign stream_matmul_16_parameter_10_data = __variable_wdata_2490;
  wire _set_flag_2221;
  assign _set_flag_2221 = matmul_16_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_2491;
  assign stream_matmul_16_source_11_data = __variable_wdata_2491;
  wire _set_flag_2222;
  assign _set_flag_2222 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2502;
  assign stream_matmul_16_parameter_12_data = __variable_wdata_2502;
  wire _set_flag_2223;
  assign _set_flag_2223 = matmul_16_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_2503;
  assign stream_matmul_16_source_13_data = __variable_wdata_2503;
  wire _set_flag_2224;
  assign _set_flag_2224 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2514;
  assign stream_matmul_16_parameter_14_data = __variable_wdata_2514;
  wire _set_flag_2225;
  assign _set_flag_2225 = matmul_16_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_2515;
  assign stream_matmul_16_source_15_data = __variable_wdata_2515;
  wire _set_flag_2226;
  assign _set_flag_2226 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2526;
  assign stream_matmul_16_parameter_16_data = __variable_wdata_2526;
  wire _set_flag_2227;
  assign _set_flag_2227 = matmul_16_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2527;
  assign stream_matmul_16_parameter_17_data = __variable_wdata_2527;
  wire _set_flag_2228;
  assign _set_flag_2228 = matmul_16_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_2528;
  assign stream_matmul_16_parameter_18_data = __variable_wdata_2528;
  wire _set_flag_2229;
  assign _set_flag_2229 = matmul_16_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_2529;
  assign stream_matmul_16_parameter_19_data = __variable_wdata_2529;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_0;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_1;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_2;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_3;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_count_0;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_count_1;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_count_2;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_count_3;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_16_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_16_source_20_pat_stride_buf_3;
  wire _set_flag_2230;
  assign _set_flag_2230 = matmul_16_comp_fsm == 3;
  assign ram_w32_l8192_id0_0_addr = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_20_source_ram_renable && (_stream_matmul_16_source_20_source_sel == 3))? _stream_matmul_16_source_20_source_ram_raddr : 
                                    (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? _stream_max_pool_serial_6_sink_6_sink_waddr : 'hx;
  assign ram_w32_l8192_id0_0_enable = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_20_source_ram_renable && (_stream_matmul_16_source_20_source_sel == 3))? 1'd1 : 
                                      (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_6_sink_wenable && (_stream_max_pool_serial_6_sink_6_sink_sel == 2))? 1'd1 : 0;
  localparam _tmp_2231 = 1;
  wire [_tmp_2231-1:0] _tmp_2232;
  assign _tmp_2232 = _stream_matmul_16_stream_oready && _stream_matmul_16_source_20_source_ram_renable && (_stream_matmul_16_source_20_source_sel == 3);
  reg [_tmp_2231-1:0] __tmp_2232_1;
  assign _stream_matmul_16_source_20_source_ram_rdata = (_stream_matmul_16_source_20_source_sel == 3)? ram_w32_l8192_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_2530;
  assign stream_matmul_16_source_20_data = __variable_wdata_2530;
  reg [32-1:0] _stream_matmul_16_source_20_source_pat_fsm_2;
  localparam _stream_matmul_16_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_matmul_16_source_20_source_pat_all_offset;
  assign _stream_matmul_16_source_20_source_pat_all_offset = _stream_matmul_16_source_20_source_offset_buf + _source_stream_matmul_16_source_20_pat_cur_offset_0 + _source_stream_matmul_16_source_20_pat_cur_offset_1 + _source_stream_matmul_16_source_20_pat_cur_offset_2 + _source_stream_matmul_16_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_0;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_1;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_2;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_3;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_count_0;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_count_1;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_count_2;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_count_3;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_16_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_16_source_21_pat_stride_buf_3;
  wire _set_flag_2233;
  assign _set_flag_2233 = matmul_16_comp_fsm == 3;
  assign ram_w32_l16384_id0_0_addr = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_21_source_ram_renable && (_stream_matmul_16_source_21_source_sel == 4))? _stream_matmul_16_source_21_source_ram_raddr : 
                                     (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? _stream_max_pool_serial_6_source_1_source_ram_raddr : 'hx;
  assign ram_w32_l16384_id0_0_enable = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_21_source_ram_renable && (_stream_matmul_16_source_21_source_sel == 4))? 1'd1 : 
                                       (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_2234 = 1;
  wire [_tmp_2234-1:0] _tmp_2235;
  assign _tmp_2235 = _stream_matmul_16_stream_oready && _stream_matmul_16_source_21_source_ram_renable && (_stream_matmul_16_source_21_source_sel == 4);
  reg [_tmp_2234-1:0] __tmp_2235_1;
  assign _stream_matmul_16_source_21_source_ram_rdata = (_stream_matmul_16_source_21_source_sel == 4)? ram_w32_l16384_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_2551;
  assign stream_matmul_16_source_21_data = __variable_wdata_2551;
  reg [32-1:0] _stream_matmul_16_source_21_source_pat_fsm_3;
  localparam _stream_matmul_16_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_matmul_16_source_21_source_pat_all_offset;
  assign _stream_matmul_16_source_21_source_pat_all_offset = _stream_matmul_16_source_21_source_offset_buf + _source_stream_matmul_16_source_21_pat_cur_offset_0 + _source_stream_matmul_16_source_21_pat_cur_offset_1 + _source_stream_matmul_16_source_21_pat_cur_offset_2 + _source_stream_matmul_16_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_0;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_1;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_2;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_3;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_count_0;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_count_1;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_count_2;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_count_3;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_16_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_16_source_22_pat_stride_buf_3;
  wire _set_flag_2236;
  assign _set_flag_2236 = matmul_16_comp_fsm == 3;
  assign ram_w32_l16384_id1_0_addr = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_22_source_ram_renable && (_stream_matmul_16_source_22_source_sel == 5))? _stream_matmul_16_source_22_source_ram_raddr : 'hx;
  assign ram_w32_l16384_id1_0_enable = (_stream_matmul_16_stream_oready && _stream_matmul_16_source_22_source_ram_renable && (_stream_matmul_16_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_2237 = 1;
  wire [_tmp_2237-1:0] _tmp_2238;
  assign _tmp_2238 = _stream_matmul_16_stream_oready && _stream_matmul_16_source_22_source_ram_renable && (_stream_matmul_16_source_22_source_sel == 5);
  reg [_tmp_2237-1:0] __tmp_2238_1;
  assign _stream_matmul_16_source_22_source_ram_rdata = (_stream_matmul_16_source_22_source_sel == 5)? ram_w32_l16384_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_2552;
  assign stream_matmul_16_source_22_data = __variable_wdata_2552;
  reg [32-1:0] _stream_matmul_16_source_22_source_pat_fsm_4;
  localparam _stream_matmul_16_source_22_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_matmul_16_source_22_source_pat_all_offset;
  assign _stream_matmul_16_source_22_source_pat_all_offset = _stream_matmul_16_source_22_source_offset_buf + _source_stream_matmul_16_source_22_pat_cur_offset_0 + _source_stream_matmul_16_source_22_pat_cur_offset_1 + _source_stream_matmul_16_source_22_pat_cur_offset_2 + _source_stream_matmul_16_source_22_pat_cur_offset_3;
  wire _set_flag_2239;
  assign _set_flag_2239 = matmul_16_comp_fsm == 3;
  reg _tmp_2240;
  reg _tmp_2241;
  reg _tmp_2242;
  reg _tmp_2243;
  reg _tmp_2244;
  reg _tmp_2245;
  reg _tmp_2246;
  reg _tmp_2247;
  reg _tmp_2248;
  reg _tmp_2249;
  reg _tmp_2250;
  reg _tmp_2251;
  reg _tmp_2252;
  reg _tmp_2253;
  reg _tmp_2254;
  reg _tmp_2255;
  reg _tmp_2256;
  reg _tmp_2257;
  reg _tmp_2258;
  reg _tmp_2259;
  reg _tmp_2260;
  reg _tmp_2261;
  reg _tmp_2262;
  reg _tmp_2263;
  reg _tmp_2264;
  reg _tmp_2265;
  reg _tmp_2266;
  reg _tmp_2267;
  reg _tmp_2268;
  reg _tmp_2269;
  reg _tmp_2270;
  reg _tmp_2271;
  reg _tmp_2272;
  reg _tmp_2273;
  localparam _tmp_2274 = 33;
  wire [_tmp_2274-1:0] _tmp_2275;
  assign _tmp_2275 = matmul_16_stream_out_local + matmul_16_out_page_comp_offset_buf;
  reg [_tmp_2274-1:0] _tmp_2276;
  reg [_tmp_2274-1:0] _tmp_2277;
  reg [_tmp_2274-1:0] _tmp_2278;
  reg [_tmp_2274-1:0] _tmp_2279;
  reg [_tmp_2274-1:0] _tmp_2280;
  reg [_tmp_2274-1:0] _tmp_2281;
  reg [_tmp_2274-1:0] _tmp_2282;
  reg [_tmp_2274-1:0] _tmp_2283;
  reg [_tmp_2274-1:0] _tmp_2284;
  reg [_tmp_2274-1:0] _tmp_2285;
  reg [_tmp_2274-1:0] _tmp_2286;
  reg [_tmp_2274-1:0] _tmp_2287;
  reg [_tmp_2274-1:0] _tmp_2288;
  reg [_tmp_2274-1:0] _tmp_2289;
  reg [_tmp_2274-1:0] _tmp_2290;
  reg [_tmp_2274-1:0] _tmp_2291;
  reg [_tmp_2274-1:0] _tmp_2292;
  reg [_tmp_2274-1:0] _tmp_2293;
  reg [_tmp_2274-1:0] _tmp_2294;
  reg [_tmp_2274-1:0] _tmp_2295;
  reg [_tmp_2274-1:0] _tmp_2296;
  reg [_tmp_2274-1:0] _tmp_2297;
  reg [_tmp_2274-1:0] _tmp_2298;
  reg [_tmp_2274-1:0] _tmp_2299;
  reg [_tmp_2274-1:0] _tmp_2300;
  reg [_tmp_2274-1:0] _tmp_2301;
  reg [_tmp_2274-1:0] _tmp_2302;
  reg [_tmp_2274-1:0] _tmp_2303;
  reg [_tmp_2274-1:0] _tmp_2304;
  reg [_tmp_2274-1:0] _tmp_2305;
  reg [_tmp_2274-1:0] _tmp_2306;
  reg [_tmp_2274-1:0] _tmp_2307;
  reg [_tmp_2274-1:0] _tmp_2308;
  reg [_tmp_2274-1:0] _tmp_2309;
  reg [32-1:0] _tmp_2310;
  reg [32-1:0] _tmp_2311;
  reg [32-1:0] _tmp_2312;
  reg [32-1:0] _tmp_2313;
  reg [32-1:0] _tmp_2314;
  reg [32-1:0] _tmp_2315;
  reg [32-1:0] _tmp_2316;
  reg [32-1:0] _tmp_2317;
  reg [32-1:0] _tmp_2318;
  reg [32-1:0] _tmp_2319;
  reg [32-1:0] _tmp_2320;
  reg [32-1:0] _tmp_2321;
  reg [32-1:0] _tmp_2322;
  reg [32-1:0] _tmp_2323;
  reg [32-1:0] _tmp_2324;
  reg [32-1:0] _tmp_2325;
  reg [32-1:0] _tmp_2326;
  reg [32-1:0] _tmp_2327;
  reg [32-1:0] _tmp_2328;
  reg [32-1:0] _tmp_2329;
  reg [32-1:0] _tmp_2330;
  reg [32-1:0] _tmp_2331;
  reg [32-1:0] _tmp_2332;
  reg [32-1:0] _tmp_2333;
  reg [32-1:0] _tmp_2334;
  reg [32-1:0] _tmp_2335;
  reg [32-1:0] _tmp_2336;
  reg [32-1:0] _tmp_2337;
  reg [32-1:0] _tmp_2338;
  reg [32-1:0] _tmp_2339;
  reg [32-1:0] _tmp_2340;
  reg [32-1:0] _tmp_2341;
  reg [32-1:0] _tmp_2342;
  reg [32-1:0] _tmp_2343;
  assign ram_w32_l128_id0_0_addr = (_stream_matmul_16_stream_oready && _stream_matmul_16_sink_33_sink_wenable && (_stream_matmul_16_sink_33_sink_sel == 6))? _stream_matmul_16_sink_33_sink_waddr : 
                                   (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? _stream_conv2d_4_source_29_source_ram_raddr : 'hx;
  assign ram_w32_l128_id0_0_wdata = (_stream_matmul_16_stream_oready && _stream_matmul_16_sink_33_sink_wenable && (_stream_matmul_16_sink_33_sink_sel == 6))? _stream_matmul_16_sink_33_sink_wdata : 'hx;
  assign ram_w32_l128_id0_0_wenable = (_stream_matmul_16_stream_oready && _stream_matmul_16_sink_33_sink_wenable && (_stream_matmul_16_sink_33_sink_sel == 6))? 1'd1 : 0;
  assign ram_w32_l128_id0_0_enable = (_stream_matmul_16_stream_oready && _stream_matmul_16_sink_33_sink_wenable && (_stream_matmul_16_sink_33_sink_sel == 6))? 1'd1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? 1'd1 : 0;
  reg [32-1:0] _stream_matmul_16_sink_33_sink_fsm_5;
  localparam _stream_matmul_16_sink_33_sink_fsm_5_init = 0;
  wire _set_flag_2344;
  assign _set_flag_2344 = matmul_16_comp_fsm == 4;
  assign _stream_matmul_16_run_flag = (_set_flag_2344)? 1 : 0;
  reg _tmp_2345;
  reg _tmp_2346;
  reg _tmp_2347;
  assign _add_tree_2_source_stop = _add_tree_2_stream_oready && 1'd0;
  reg _tmp_2348;
  reg _tmp_2349;
  reg _tmp_2350;
  assign _add_tree_2_sink_start = _tmp_2350;
  reg _tmp_2351;
  reg _tmp_2352;
  reg _tmp_2353;
  assign _add_tree_2_sink_stop = _tmp_2353;
  reg _tmp_2354;
  reg _tmp_2355;
  reg _tmp_2356;
  assign _add_tree_2_sink_busy = _tmp_2356;
  reg _tmp_2357;
  assign _add_tree_2_busy = _add_tree_2_source_busy || _add_tree_2_sink_busy || _add_tree_2_busy_reg;
  reg _tmp_2358;
  reg _tmp_2359;
  reg _tmp_2360;
  assign _add_tree_3_source_stop = _add_tree_3_stream_oready && 1'd0;
  reg _tmp_2361;
  reg _tmp_2362;
  reg _tmp_2363;
  assign _add_tree_3_sink_start = _tmp_2363;
  reg _tmp_2364;
  reg _tmp_2365;
  reg _tmp_2366;
  assign _add_tree_3_sink_stop = _tmp_2366;
  reg _tmp_2367;
  reg _tmp_2368;
  reg _tmp_2369;
  assign _add_tree_3_sink_busy = _tmp_2369;
  reg _tmp_2370;
  assign _add_tree_3_busy = _add_tree_3_source_busy || _add_tree_3_sink_busy || _add_tree_3_busy_reg;
  reg _tmp_2371;
  reg _tmp_2372;
  reg _tmp_2373;
  reg _tmp_2374;
  reg _tmp_2375;
  reg _tmp_2376;
  reg [1-1:0] __variable_wdata_2450;
  assign stream_matmul_16__reduce_reset_data = __variable_wdata_2450;
  reg _tmp_2377;
  reg _tmp_2378;
  reg _tmp_2379;
  reg _tmp_2380;
  assign _stream_matmul_16_source_stop = _stream_matmul_16_stream_oready && (_stream_matmul_16_source_11_idle && _stream_matmul_16_source_13_idle && _stream_matmul_16_source_15_idle && _stream_matmul_16_source_20_idle && _stream_matmul_16_source_21_idle && _stream_matmul_16_source_22_idle && _stream_matmul_16_source_7_idle && _stream_matmul_16_source_9_idle && (_stream_matmul_16_fsm == 3));
  localparam _tmp_2381 = 1;
  wire [_tmp_2381-1:0] _tmp_2382;
  assign _tmp_2382 = _stream_matmul_16_source_11_idle && _stream_matmul_16_source_13_idle && _stream_matmul_16_source_15_idle && _stream_matmul_16_source_20_idle && _stream_matmul_16_source_21_idle && _stream_matmul_16_source_22_idle && _stream_matmul_16_source_7_idle && _stream_matmul_16_source_9_idle && (_stream_matmul_16_fsm == 3);
  reg [_tmp_2381-1:0] _tmp_2383;
  localparam _tmp_2384 = 1;
  wire [_tmp_2384-1:0] _tmp_2385;
  assign _tmp_2385 = _stream_matmul_16_source_11_idle && _stream_matmul_16_source_13_idle && _stream_matmul_16_source_15_idle && _stream_matmul_16_source_20_idle && _stream_matmul_16_source_21_idle && _stream_matmul_16_source_22_idle && _stream_matmul_16_source_7_idle && _stream_matmul_16_source_9_idle && (_stream_matmul_16_fsm == 3);
  reg [_tmp_2384-1:0] _tmp_2386;
  reg _tmp_2387;
  reg _tmp_2388;
  reg _tmp_2389;
  reg _tmp_2390;
  reg _tmp_2391;
  reg _tmp_2392;
  reg _tmp_2393;
  reg _tmp_2394;
  reg _tmp_2395;
  reg _tmp_2396;
  reg _tmp_2397;
  reg _tmp_2398;
  reg _tmp_2399;
  reg _tmp_2400;
  reg _tmp_2401;
  reg _tmp_2402;
  reg _tmp_2403;
  reg _tmp_2404;
  reg _tmp_2405;
  reg _tmp_2406;
  reg _tmp_2407;
  reg _tmp_2408;
  reg _tmp_2409;
  reg _tmp_2410;
  reg _tmp_2411;
  reg _tmp_2412;
  reg _tmp_2413;
  reg _tmp_2414;
  reg _tmp_2415;
  reg _tmp_2416;
  reg _tmp_2417;
  reg _tmp_2418;
  reg _tmp_2419;
  reg _tmp_2420;
  assign _stream_matmul_16_sink_start = _tmp_2420;
  reg _tmp_2421;
  reg _tmp_2422;
  reg _tmp_2423;
  reg _tmp_2424;
  reg _tmp_2425;
  reg _tmp_2426;
  reg _tmp_2427;
  reg _tmp_2428;
  reg _tmp_2429;
  reg _tmp_2430;
  reg _tmp_2431;
  reg _tmp_2432;
  reg _tmp_2433;
  reg _tmp_2434;
  reg _tmp_2435;
  reg _tmp_2436;
  reg _tmp_2437;
  reg _tmp_2438;
  reg _tmp_2439;
  reg _tmp_2440;
  reg _tmp_2441;
  reg _tmp_2442;
  reg _tmp_2443;
  reg _tmp_2444;
  reg _tmp_2445;
  reg _tmp_2446;
  reg _tmp_2447;
  reg _tmp_2448;
  reg _tmp_2449;
  reg _tmp_2450;
  reg _tmp_2451;
  reg _tmp_2452;
  reg _tmp_2453;
  reg _tmp_2454;
  assign _stream_matmul_16_sink_stop = _tmp_2454;
  reg _tmp_2455;
  reg _tmp_2456;
  reg _tmp_2457;
  reg _tmp_2458;
  reg _tmp_2459;
  reg _tmp_2460;
  reg _tmp_2461;
  reg _tmp_2462;
  reg _tmp_2463;
  reg _tmp_2464;
  reg _tmp_2465;
  reg _tmp_2466;
  reg _tmp_2467;
  reg _tmp_2468;
  reg _tmp_2469;
  reg _tmp_2470;
  reg _tmp_2471;
  reg _tmp_2472;
  reg _tmp_2473;
  reg _tmp_2474;
  reg _tmp_2475;
  reg _tmp_2476;
  reg _tmp_2477;
  reg _tmp_2478;
  reg _tmp_2479;
  reg _tmp_2480;
  reg _tmp_2481;
  reg _tmp_2482;
  reg _tmp_2483;
  reg _tmp_2484;
  reg _tmp_2485;
  reg _tmp_2486;
  reg _tmp_2487;
  reg _tmp_2488;
  assign _stream_matmul_16_sink_busy = _tmp_2488;
  reg _tmp_2489;
  assign _stream_matmul_16_busy = _stream_matmul_16_source_busy || _stream_matmul_16_sink_busy || _stream_matmul_16_busy_reg;
  wire matmul_16_dma_out_mask_0;
  assign matmul_16_dma_out_mask_0 = matmul_16_out_row_count + 0 >= cparam_matmul_16_out_num_row;
  wire [32-1:0] mask_addr_shifted_2490;
  assign mask_addr_shifted_2490 = matmul_16_objaddr + (matmul_16_out_base_offset + cparam_matmul_16_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_2491;
  assign mask_addr_masked_2491 = mask_addr_shifted_2490 << 2;
  reg [32-1:0] read_burst_fsm_42;
  localparam read_burst_fsm_42_init = 0;
  reg [7-1:0] read_burst_addr_2492;
  reg [7-1:0] read_burst_stride_2493;
  reg [33-1:0] read_burst_length_2494;
  reg read_burst_rvalid_2495;
  reg read_burst_rlast_2496;
  assign ram_w32_l128_id0_1_addr = ((read_burst_fsm_42 == 1) && (!read_burst_rvalid_2495 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_2492 : 
                                   ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? write_burst_addr_90 : 'hx;
  assign ram_w32_l128_id0_1_enable = ((read_burst_fsm_42 == 1) && (!read_burst_rvalid_2495 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                     ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? 1'd1 : 0;
  localparam _tmp_2497 = 1;
  wire [_tmp_2497-1:0] _tmp_2498;
  assign _tmp_2498 = (read_burst_fsm_42 == 1) && (!read_burst_rvalid_2495 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_2497-1:0] __tmp_2498_1;
  wire [32-1:0] read_burst_rdata_2499;
  assign read_burst_rdata_2499 = ram_w32_l128_id0_1_rdata;
  assign _maxi_write_req_fifo_deq = ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) && !_maxi_write_req_fifo_empty)? 1 : 0;
  reg _maxi_wdata_cond_2_1;
  wire matmul_16_update_filter;
  assign matmul_16_update_filter = (cparam_matmul_16_data_stationary == 0) && (matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count) || (cparam_matmul_16_data_stationary == 1) && !cparam_matmul_16_keep_filter;
  wire matmul_16_update_act;
  assign matmul_16_update_act = (cparam_matmul_16_data_stationary == 1) && (matmul_16_och_count >= cparam_matmul_16_max_och_count) || (cparam_matmul_16_data_stationary == 0);
  wire matmul_16_mux_next_dma_flag_0;
  assign matmul_16_mux_next_dma_flag_0 = (matmul_16_row_select == 0)? (matmul_16_row_count >= cparam_matmul_16_max_row_count)? 1 : cparam_matmul_16_dma_flag_conds_0 : 1'd0;

  always @(posedge CLK) begin
    _RESETN_inv_1 <= RESETN_inv;
    _RESETN_inv_2 <= _RESETN_inv_1;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_awaddr <= 0;
      maxi_awlen <= 0;
      maxi_awvalid <= 0;
      _maxi_waddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_waddr_cond_0_1) begin
        maxi_awvalid <= 0;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid))) begin
        maxi_awaddr <= _maxi_write_global_addr;
        maxi_awlen <= _maxi_write_cur_global_size - 1;
        maxi_awvalid <= 1;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid)) && (_maxi_write_cur_global_size == 0)) begin
        maxi_awvalid <= 0;
      end 
      _maxi_waddr_cond_0_1 <= 1;
      if(maxi_awvalid && !maxi_awready) begin
        maxi_awvalid <= maxi_awvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_wdata_sb_0 <= 0;
      _maxi_wvalid_sb_0 <= 0;
      _maxi_wlast_sb_0 <= 0;
      _maxi_wstrb_sb_0 <= 0;
      _maxi_wdata_cond_0_1 <= 0;
      _maxi_wdata_cond_1_1 <= 0;
      _maxi_wdata_cond_2_1 <= 0;
    end else begin
      if(_maxi_wdata_cond_0_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_1_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_2_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_2040 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_2044;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_2041 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_0_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_2166 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_2170;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_2167 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_1_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_2495 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_2499;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_2496 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_2_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_writedata_data_6 <= 0;
      _sb_maxi_writedata_valid_7 <= 0;
      _sb_maxi_writedata_tmp_data_9 <= 0;
      _sb_maxi_writedata_tmp_valid_10 <= 0;
    end else begin
      if(_sb_maxi_writedata_m_ready_5 || !_sb_maxi_writedata_valid_7) begin
        _sb_maxi_writedata_data_6 <= _sb_maxi_writedata_next_data_11;
        _sb_maxi_writedata_valid_7 <= _sb_maxi_writedata_next_valid_12;
      end 
      if(!_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_valid_7 && !_sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_data_9 <= _sb_maxi_writedata_s_data_3;
        _sb_maxi_writedata_tmp_valid_10 <= _sb_maxi_writedata_s_valid_4;
      end 
      if(_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_valid_10 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_araddr <= 0;
      maxi_arlen <= 0;
      maxi_arvalid <= 0;
      _maxi_raddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_raddr_cond_0_1) begin
        maxi_arvalid <= 0;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        maxi_araddr <= _maxi_read_global_addr;
        maxi_arlen <= _maxi_read_cur_global_size - 1;
        maxi_arvalid <= 1;
      end 
      _maxi_raddr_cond_0_1 <= 1;
      if(maxi_arvalid && !maxi_arready) begin
        maxi_arvalid <= maxi_arvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_readdata_data_21 <= 0;
      _sb_maxi_readdata_valid_22 <= 0;
      _sb_maxi_readdata_tmp_data_24 <= 0;
      _sb_maxi_readdata_tmp_valid_25 <= 0;
    end else begin
      if(_sb_maxi_readdata_m_ready_20 || !_sb_maxi_readdata_valid_22) begin
        _sb_maxi_readdata_data_21 <= _sb_maxi_readdata_next_data_26;
        _sb_maxi_readdata_valid_22 <= _sb_maxi_readdata_next_valid_27;
      end 
      if(!_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_valid_22 && !_sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_data_24 <= _sb_maxi_readdata_s_data_18;
        _sb_maxi_readdata_tmp_valid_25 <= _sb_maxi_readdata_s_valid_19;
      end 
      if(_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_valid_25 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_outstanding_wcount <= 0;
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= 0;
      _maxi_read_op_sel <= 0;
      _maxi_read_global_addr <= 0;
      _maxi_read_global_size <= 0;
      _maxi_read_local_addr <= 0;
      _maxi_read_local_stride <= 0;
      _maxi_read_local_size <= 0;
      _maxi_read_local_blocksize <= 0;
      _maxi_read_req_busy <= 0;
      _maxi_read_cur_global_size <= 0;
      _maxi_read_data_busy <= 0;
      _maxi_read_op_sel_buf <= 0;
      _maxi_read_local_addr_buf <= 0;
      _maxi_read_local_stride_buf <= 0;
      _maxi_read_local_size_buf <= 0;
      _maxi_read_local_blocksize_buf <= 0;
      _maxi_write_op_sel <= 0;
      _maxi_write_global_addr <= 0;
      _maxi_write_global_size <= 0;
      _maxi_write_local_addr <= 0;
      _maxi_write_local_stride <= 0;
      _maxi_write_local_size <= 0;
      _maxi_write_local_blocksize <= 0;
      _maxi_write_req_busy <= 0;
      _maxi_write_cur_global_size <= 0;
      _maxi_write_data_busy <= 0;
      _maxi_write_op_sel_buf <= 0;
      _maxi_write_local_addr_buf <= 0;
      _maxi_write_local_stride_buf <= 0;
      _maxi_write_size_buf <= 0;
      _maxi_write_local_blocksize_buf <= 0;
    end else begin
      if(maxi_awvalid && maxi_awready && !(maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount < 7)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount + 1;
      end 
      if(!(maxi_awvalid && maxi_awready) && (maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount > 0)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount - 1;
      end 
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= _saxi_register_32;
      if((control_conv2d_4 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 1;
        _maxi_read_global_addr <= mask_addr_masked_55;
        _maxi_read_global_size <= cparam_conv2d_4_bias_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_4_bias_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && _maxi_read_start) begin
        _maxi_read_req_busy <= 1;
      end 
      if(_maxi_read_start && _maxi_read_req_fifo_almost_full) begin
        _maxi_read_start <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256) && ((mask_addr_masked_65 & 4095) + (_maxi_read_global_size << 2) >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_67 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_69 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256)) begin
        _maxi_read_cur_global_size <= _maxi_read_global_size;
        _maxi_read_global_size <= 0;
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && ((mask_addr_masked_71 & 4095) + 1024 >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_73 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_75 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
        _maxi_read_cur_global_size <= 256;
        _maxi_read_global_size <= _maxi_read_global_size - 256;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        _maxi_read_global_addr <= _maxi_read_global_addr + (_maxi_read_cur_global_size << 2);
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
        _maxi_read_req_busy <= 0;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 2;
        _maxi_read_global_addr <= mask_addr_masked_81;
        _maxi_read_global_size <= cparam_conv2d_4_scale_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_4_scale_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 3;
        _maxi_read_global_addr <= mask_addr_masked_87;
        _maxi_read_global_size <= cparam_conv2d_4_filter_read_size;
        _maxi_read_local_addr <= conv2d_4_filter_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_4_filter_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_4_filter_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 4;
        _maxi_read_global_addr <= mask_addr_masked_201;
        _maxi_read_global_size <= cparam_conv2d_4_act_read_size;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_4_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_4_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 17) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 5;
        _maxi_read_global_addr <= mask_addr_masked_225;
        _maxi_read_global_size <= cparam_conv2d_4_act_read_size;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_1;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_4_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_4_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 20) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 6;
        _maxi_read_global_addr <= mask_addr_masked_249;
        _maxi_read_global_size <= cparam_conv2d_4_act_read_size;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_2;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_4_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_4_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 29) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_2008;
        _maxi_write_global_size <= conv2d_4_next_out_write_size;
        _maxi_write_local_addr <= conv2d_4_out_laddr_offset + conv2d_4_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= conv2d_4_next_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && _maxi_write_start) begin
        _maxi_write_req_busy <= 1;
      end 
      if(_maxi_write_start && _maxi_write_req_fifo_almost_full) begin
        _maxi_write_start <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256) && ((mask_addr_masked_2018 & 4095) + (_maxi_write_global_size << 2) >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_2020 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_2022 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256)) begin
        _maxi_write_cur_global_size <= _maxi_write_global_size;
        _maxi_write_global_size <= 0;
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && ((mask_addr_masked_2024 & 4095) + 1024 >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_2026 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_2028 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
        _maxi_write_cur_global_size <= 256;
        _maxi_write_global_size <= _maxi_write_global_size - 256;
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))) begin
        _maxi_write_global_addr <= _maxi_write_global_addr + (_maxi_write_cur_global_size << 2);
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) && (_maxi_write_global_size == 0)) begin
        _maxi_write_req_busy <= 0;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_2040 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_2040 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_2041) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_max_pool_serial_6 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_2046;
        _maxi_read_global_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_addr <= max_pool_serial_6_act_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_max_pool_serial_6 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_2052;
        _maxi_read_global_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_addr <= max_pool_serial_6_act_page_dma_offset + cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_max_pool_serial_6 == 15) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 2;
        _maxi_write_global_addr <= mask_addr_masked_2162;
        _maxi_write_global_size <= cparam_max_pool_serial_6_out_write_size;
        _maxi_write_local_addr <= max_pool_serial_6_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= cparam_max_pool_serial_6_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_2166 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_2166 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_2167) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_matmul_16 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 8;
        _maxi_read_global_addr <= mask_addr_masked_2172;
        _maxi_read_global_size <= cparam_matmul_16_bias_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_16_bias_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_16 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 9;
        _maxi_read_global_addr <= mask_addr_masked_2178;
        _maxi_read_global_size <= cparam_matmul_16_scale_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_16_scale_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_16 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 10;
        _maxi_read_global_addr <= mask_addr_masked_2184;
        _maxi_read_global_size <= cparam_matmul_16_filter_read_size;
        _maxi_read_local_addr <= matmul_16_filter_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_16_filter_read_size;
        _maxi_read_local_blocksize <= cparam_matmul_16_filter_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_16 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 11;
        _maxi_read_global_addr <= mask_addr_masked_2202;
        _maxi_read_global_size <= cparam_matmul_16_act_read_size;
        _maxi_read_local_addr <= matmul_16_act_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_16_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 11))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_16 == 23) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 3;
        _maxi_write_global_addr <= mask_addr_masked_2491;
        _maxi_write_global_size <= matmul_16_next_out_write_size;
        _maxi_write_local_addr <= matmul_16_out_laddr_offset + matmul_16_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= matmul_16_next_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_2495 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_2495 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_2496) begin
        _maxi_write_data_busy <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_read_req_fifo <= 0;
      __tmp_63_1 <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full && (_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty)) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo;
      end else if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo + 1;
      end else if(_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo - 1;
      end 
      __tmp_63_1 <= _tmp_63;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_write_req_fifo <= 0;
      __tmp_2016_1 <= 0;
      __tmp_2036_1 <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full && (_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty)) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo;
      end else if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo + 1;
      end else if(_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo - 1;
      end 
      __tmp_2016_1 <= _tmp_2016;
      __tmp_2036_1 <= _tmp_2036;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_rdata <= 0;
      saxi_rvalid <= 0;
      _saxi_rdata_cond_0_1 <= 0;
    end else begin
      if(_saxi_rdata_cond_0_1) begin
        saxi_rvalid <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid)) begin
        saxi_rdata <= axislite_rdata_46;
        saxi_rvalid <= 1;
      end 
      _saxi_rdata_cond_0_1 <= 1;
      if(saxi_rvalid && !saxi_rready) begin
        saxi_rvalid <= saxi_rvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_bvalid <= 0;
      prev_awvalid_43 <= 0;
      prev_arvalid_44 <= 0;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      addr_40 <= 0;
      _saxi_register_0 <= 0;
      _saxi_flag_0 <= 0;
      _saxi_register_1 <= 0;
      _saxi_flag_1 <= 0;
      _saxi_register_2 <= 0;
      _saxi_flag_2 <= 0;
      _saxi_register_3 <= 0;
      _saxi_flag_3 <= 0;
      _saxi_register_4 <= 0;
      _saxi_flag_4 <= 0;
      _saxi_register_5 <= 0;
      _saxi_flag_5 <= 0;
      _saxi_register_6 <= 0;
      _saxi_flag_6 <= 0;
      _saxi_register_7 <= 0;
      _saxi_flag_7 <= 0;
      _saxi_register_8 <= 0;
      _saxi_flag_8 <= 0;
      _saxi_register_9 <= 0;
      _saxi_flag_9 <= 0;
      _saxi_register_10 <= 0;
      _saxi_flag_10 <= 0;
      _saxi_register_11 <= 0;
      _saxi_flag_11 <= 0;
      _saxi_register_12 <= 0;
      _saxi_flag_12 <= 0;
      _saxi_register_13 <= 0;
      _saxi_flag_13 <= 0;
      _saxi_register_14 <= 0;
      _saxi_flag_14 <= 0;
      _saxi_register_15 <= 0;
      _saxi_flag_15 <= 0;
      _saxi_register_16 <= 0;
      _saxi_flag_16 <= 0;
      _saxi_register_17 <= 0;
      _saxi_flag_17 <= 0;
      _saxi_register_18 <= 0;
      _saxi_flag_18 <= 0;
      _saxi_register_19 <= 0;
      _saxi_flag_19 <= 0;
      _saxi_register_20 <= 0;
      _saxi_flag_20 <= 0;
      _saxi_register_21 <= 0;
      _saxi_flag_21 <= 0;
      _saxi_register_22 <= 0;
      _saxi_flag_22 <= 0;
      _saxi_register_23 <= 0;
      _saxi_flag_23 <= 0;
      _saxi_register_24 <= 0;
      _saxi_flag_24 <= 0;
      _saxi_register_25 <= 0;
      _saxi_flag_25 <= 0;
      _saxi_register_26 <= 0;
      _saxi_flag_26 <= 0;
      _saxi_register_27 <= 0;
      _saxi_flag_27 <= 0;
      _saxi_register_28 <= 0;
      _saxi_flag_28 <= 0;
      _saxi_register_29 <= 0;
      _saxi_flag_29 <= 0;
      _saxi_register_30 <= 0;
      _saxi_flag_30 <= 0;
      _saxi_register_31 <= 8679104;
      _saxi_flag_31 <= 0;
      _saxi_register_32 <= 0;
      _saxi_flag_32 <= 0;
      _saxi_register_33 <= 8481984;
      _saxi_flag_33 <= 0;
      _saxi_register_34 <= 0;
      _saxi_flag_34 <= 0;
      _saxi_register_35 <= 64;
      _saxi_flag_35 <= 0;
      _saxi_register_36 <= 8256;
      _saxi_flag_36 <= 0;
      _saxi_register_11[0] <= (0 >> 0) & 1'd1;
      _saxi_register_9[0] <= (0 >> 0) & 1'd1;
      _saxi_register_11[1] <= (0 >> 1) & 1'd1;
      _saxi_register_9[1] <= (0 >> 1) & 1'd1;
      _saxi_register_11[2] <= (0 >> 2) & 1'd1;
      _saxi_register_9[2] <= (0 >> 2) & 1'd1;
      _saxi_register_11[3] <= (0 >> 3) & 1'd1;
      _saxi_register_9[3] <= (0 >> 3) & 1'd1;
      _saxi_register_11[4] <= (0 >> 4) & 1'd1;
      _saxi_register_9[4] <= (0 >> 4) & 1'd1;
      _saxi_register_11[5] <= (0 >> 5) & 1'd1;
      _saxi_register_9[5] <= (0 >> 5) & 1'd1;
      _saxi_register_11[6] <= (0 >> 6) & 1'd1;
      _saxi_register_9[6] <= (0 >> 6) & 1'd1;
      _saxi_register_11[7] <= (0 >> 7) & 1'd1;
      _saxi_register_9[7] <= (0 >> 7) & 1'd1;
      _saxi_register_11[8] <= (0 >> 8) & 1'd1;
      _saxi_register_9[8] <= (0 >> 8) & 1'd1;
      _saxi_register_11[9] <= (0 >> 9) & 1'd1;
      _saxi_register_9[9] <= (0 >> 9) & 1'd1;
      _saxi_register_11[10] <= (0 >> 10) & 1'd1;
      _saxi_register_9[10] <= (0 >> 10) & 1'd1;
      _saxi_register_11[11] <= (0 >> 11) & 1'd1;
      _saxi_register_9[11] <= (0 >> 11) & 1'd1;
      _saxi_register_11[12] <= (0 >> 12) & 1'd1;
      _saxi_register_9[12] <= (0 >> 12) & 1'd1;
      _saxi_register_11[13] <= (0 >> 13) & 1'd1;
      _saxi_register_9[13] <= (0 >> 13) & 1'd1;
      _saxi_register_11[14] <= (0 >> 14) & 1'd1;
      _saxi_register_9[14] <= (0 >> 14) & 1'd1;
      _saxi_register_11[15] <= (0 >> 15) & 1'd1;
      _saxi_register_9[15] <= (0 >> 15) & 1'd1;
      _saxi_register_11[16] <= (0 >> 16) & 1'd1;
      _saxi_register_9[16] <= (0 >> 16) & 1'd1;
      _saxi_register_11[17] <= (0 >> 17) & 1'd1;
      _saxi_register_9[17] <= (0 >> 17) & 1'd1;
      _saxi_register_11[18] <= (0 >> 18) & 1'd1;
      _saxi_register_9[18] <= (0 >> 18) & 1'd1;
      _saxi_register_11[19] <= (0 >> 19) & 1'd1;
      _saxi_register_9[19] <= (0 >> 19) & 1'd1;
      _saxi_register_11[20] <= (0 >> 20) & 1'd1;
      _saxi_register_9[20] <= (0 >> 20) & 1'd1;
      _saxi_register_11[21] <= (0 >> 21) & 1'd1;
      _saxi_register_9[21] <= (0 >> 21) & 1'd1;
      _saxi_register_11[22] <= (0 >> 22) & 1'd1;
      _saxi_register_9[22] <= (0 >> 22) & 1'd1;
      _saxi_register_11[23] <= (0 >> 23) & 1'd1;
      _saxi_register_9[23] <= (0 >> 23) & 1'd1;
      _saxi_register_11[24] <= (0 >> 24) & 1'd1;
      _saxi_register_9[24] <= (0 >> 24) & 1'd1;
      _saxi_register_11[25] <= (0 >> 25) & 1'd1;
      _saxi_register_9[25] <= (0 >> 25) & 1'd1;
      _saxi_register_11[26] <= (0 >> 26) & 1'd1;
      _saxi_register_9[26] <= (0 >> 26) & 1'd1;
      _saxi_register_11[27] <= (0 >> 27) & 1'd1;
      _saxi_register_9[27] <= (0 >> 27) & 1'd1;
      _saxi_register_11[28] <= (0 >> 28) & 1'd1;
      _saxi_register_9[28] <= (0 >> 28) & 1'd1;
      _saxi_register_11[29] <= (0 >> 29) & 1'd1;
      _saxi_register_9[29] <= (0 >> 29) & 1'd1;
      _saxi_register_11[30] <= (0 >> 30) & 1'd1;
      _saxi_register_9[30] <= (0 >> 30) & 1'd1;
      _saxi_register_11[31] <= (0 >> 31) & 1'd1;
      _saxi_register_9[31] <= (0 >> 31) & 1'd1;
      internal_state_counter <= 0;
    end else begin
      if(saxi_bvalid && saxi_bready) begin
        saxi_bvalid <= 0;
      end 
      if(saxi_wvalid && saxi_wready) begin
        saxi_bvalid <= 1;
      end 
      prev_awvalid_43 <= saxi_awvalid;
      prev_arvalid_44 <= saxi_arvalid;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      if(saxi_awready && saxi_awvalid && !saxi_bvalid) begin
        addr_40 <= saxi_awaddr;
        writevalid_41 <= 1;
      end else if(saxi_arready && saxi_arvalid) begin
        addr_40 <= saxi_araddr;
        readvalid_42 <= 1;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= axislite_resetval_48;
        _saxi_flag_0 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= axislite_resetval_48;
        _saxi_flag_1 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= axislite_resetval_48;
        _saxi_flag_2 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= axislite_resetval_48;
        _saxi_flag_3 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= axislite_resetval_48;
        _saxi_flag_4 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= axislite_resetval_48;
        _saxi_flag_5 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= axislite_resetval_48;
        _saxi_flag_6 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= axislite_resetval_48;
        _saxi_flag_7 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= axislite_resetval_48;
        _saxi_flag_8 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= axislite_resetval_48;
        _saxi_flag_9 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= axislite_resetval_48;
        _saxi_flag_10 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= axislite_resetval_48;
        _saxi_flag_11 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= axislite_resetval_48;
        _saxi_flag_12 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= axislite_resetval_48;
        _saxi_flag_13 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= axislite_resetval_48;
        _saxi_flag_14 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= axislite_resetval_48;
        _saxi_flag_15 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= axislite_resetval_48;
        _saxi_flag_16 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= axislite_resetval_48;
        _saxi_flag_17 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= axislite_resetval_48;
        _saxi_flag_18 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= axislite_resetval_48;
        _saxi_flag_19 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= axislite_resetval_48;
        _saxi_flag_20 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= axislite_resetval_48;
        _saxi_flag_21 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= axislite_resetval_48;
        _saxi_flag_22 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= axislite_resetval_48;
        _saxi_flag_23 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= axislite_resetval_48;
        _saxi_flag_24 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= axislite_resetval_48;
        _saxi_flag_25 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= axislite_resetval_48;
        _saxi_flag_26 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= axislite_resetval_48;
        _saxi_flag_27 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= axislite_resetval_48;
        _saxi_flag_28 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= axislite_resetval_48;
        _saxi_flag_29 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= axislite_resetval_48;
        _saxi_flag_30 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= axislite_resetval_48;
        _saxi_flag_31 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= axislite_resetval_48;
        _saxi_flag_32 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= axislite_resetval_48;
        _saxi_flag_33 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= axislite_resetval_48;
        _saxi_flag_34 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= axislite_resetval_48;
        _saxi_flag_35 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= axislite_resetval_48;
        _saxi_flag_36 <= 0;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= saxi_wdata;
      end 
      if(_saxi_register_11[0] == 1) begin
        _saxi_register_11[0] <= 0;
        _saxi_register_9[0] <= 0;
      end 
      if(_saxi_register_11[1] == 1) begin
        _saxi_register_11[1] <= 0;
        _saxi_register_9[1] <= 0;
      end 
      if(_saxi_register_11[2] == 1) begin
        _saxi_register_11[2] <= 0;
        _saxi_register_9[2] <= 0;
      end 
      if(_saxi_register_11[3] == 1) begin
        _saxi_register_11[3] <= 0;
        _saxi_register_9[3] <= 0;
      end 
      if(_saxi_register_11[4] == 1) begin
        _saxi_register_11[4] <= 0;
        _saxi_register_9[4] <= 0;
      end 
      if(_saxi_register_11[5] == 1) begin
        _saxi_register_11[5] <= 0;
        _saxi_register_9[5] <= 0;
      end 
      if(_saxi_register_11[6] == 1) begin
        _saxi_register_11[6] <= 0;
        _saxi_register_9[6] <= 0;
      end 
      if(_saxi_register_11[7] == 1) begin
        _saxi_register_11[7] <= 0;
        _saxi_register_9[7] <= 0;
      end 
      if(_saxi_register_11[8] == 1) begin
        _saxi_register_11[8] <= 0;
        _saxi_register_9[8] <= 0;
      end 
      if(_saxi_register_11[9] == 1) begin
        _saxi_register_11[9] <= 0;
        _saxi_register_9[9] <= 0;
      end 
      if(_saxi_register_11[10] == 1) begin
        _saxi_register_11[10] <= 0;
        _saxi_register_9[10] <= 0;
      end 
      if(_saxi_register_11[11] == 1) begin
        _saxi_register_11[11] <= 0;
        _saxi_register_9[11] <= 0;
      end 
      if(_saxi_register_11[12] == 1) begin
        _saxi_register_11[12] <= 0;
        _saxi_register_9[12] <= 0;
      end 
      if(_saxi_register_11[13] == 1) begin
        _saxi_register_11[13] <= 0;
        _saxi_register_9[13] <= 0;
      end 
      if(_saxi_register_11[14] == 1) begin
        _saxi_register_11[14] <= 0;
        _saxi_register_9[14] <= 0;
      end 
      if(_saxi_register_11[15] == 1) begin
        _saxi_register_11[15] <= 0;
        _saxi_register_9[15] <= 0;
      end 
      if(_saxi_register_11[16] == 1) begin
        _saxi_register_11[16] <= 0;
        _saxi_register_9[16] <= 0;
      end 
      if(_saxi_register_11[17] == 1) begin
        _saxi_register_11[17] <= 0;
        _saxi_register_9[17] <= 0;
      end 
      if(_saxi_register_11[18] == 1) begin
        _saxi_register_11[18] <= 0;
        _saxi_register_9[18] <= 0;
      end 
      if(_saxi_register_11[19] == 1) begin
        _saxi_register_11[19] <= 0;
        _saxi_register_9[19] <= 0;
      end 
      if(_saxi_register_11[20] == 1) begin
        _saxi_register_11[20] <= 0;
        _saxi_register_9[20] <= 0;
      end 
      if(_saxi_register_11[21] == 1) begin
        _saxi_register_11[21] <= 0;
        _saxi_register_9[21] <= 0;
      end 
      if(_saxi_register_11[22] == 1) begin
        _saxi_register_11[22] <= 0;
        _saxi_register_9[22] <= 0;
      end 
      if(_saxi_register_11[23] == 1) begin
        _saxi_register_11[23] <= 0;
        _saxi_register_9[23] <= 0;
      end 
      if(_saxi_register_11[24] == 1) begin
        _saxi_register_11[24] <= 0;
        _saxi_register_9[24] <= 0;
      end 
      if(_saxi_register_11[25] == 1) begin
        _saxi_register_11[25] <= 0;
        _saxi_register_9[25] <= 0;
      end 
      if(_saxi_register_11[26] == 1) begin
        _saxi_register_11[26] <= 0;
        _saxi_register_9[26] <= 0;
      end 
      if(_saxi_register_11[27] == 1) begin
        _saxi_register_11[27] <= 0;
        _saxi_register_9[27] <= 0;
      end 
      if(_saxi_register_11[28] == 1) begin
        _saxi_register_11[28] <= 0;
        _saxi_register_9[28] <= 0;
      end 
      if(_saxi_register_11[29] == 1) begin
        _saxi_register_11[29] <= 0;
        _saxi_register_9[29] <= 0;
      end 
      if(_saxi_register_11[30] == 1) begin
        _saxi_register_11[30] <= 0;
        _saxi_register_9[30] <= 0;
      end 
      if(_saxi_register_11[31] == 1) begin
        _saxi_register_11[31] <= 0;
        _saxi_register_9[31] <= 0;
      end 
      if(irq_busy_edge_51) begin
        _saxi_register_9[0] <= irq_busy_edge_51;
      end 
      if(irq_extern_edge_53) begin
        _saxi_register_9[1] <= irq_extern_edge_53;
      end 
      if(main_fsm == 0) begin
        _saxi_register_5 <= 0;
        _saxi_register_6 <= 0;
        _saxi_register_7 <= 0;
      end 
      if(main_fsm == 1) begin
        internal_state_counter <= 0;
        _saxi_register_12 <= 0;
      end else if(main_fsm == _saxi_register_13) begin
        if(internal_state_counter == _saxi_register_14) begin
          internal_state_counter <= 0;
          _saxi_register_12 <= _saxi_register_12 + 1;
        end else begin
          internal_state_counter <= internal_state_counter + 1;
        end
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_0 <= 1;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_1 <= 1;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_2 <= 1;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_3 <= 1;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_4 <= 1;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 1) && 1) begin
        _saxi_register_5 <= 1;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_6 <= 1;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_7 <= 1;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_8 <= 1;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_9 <= 1;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_10 <= 1;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_11 <= 1;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_12 <= 1;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_13 <= 1;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_14 <= 1;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_15 <= 1;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_16 <= 1;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_17 <= 1;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_18 <= 1;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_19 <= 1;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_20 <= 1;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_21 <= 1;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_22 <= 1;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_23 <= 1;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_24 <= 1;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_25 <= 1;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_26 <= 1;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_27 <= 1;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_28 <= 1;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_29 <= 1;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_30 <= 1;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_31 <= 1;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_32 <= 1;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_33 <= 1;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_34 <= 1;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_35 <= 1;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_36 <= 1;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 2) && 1) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 54) && 1) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 54) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
    end
  end

  localparam _saxi_register_fsm_1 = 1;
  localparam _saxi_register_fsm_2 = 2;
  localparam _saxi_register_fsm_3 = 3;
  localparam _saxi_register_fsm_4 = 4;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _saxi_register_fsm <= _saxi_register_fsm_init;
      axis_maskaddr_45 <= 0;
    end else begin
      case(_saxi_register_fsm)
        _saxi_register_fsm_init: begin
          if(readvalid_42 || writevalid_41) begin
            axis_maskaddr_45 <= (addr_40 >> _saxi_shift) & _saxi_mask;
          end 
          if(readvalid_42) begin
            _saxi_register_fsm <= _saxi_register_fsm_1;
          end 
          if(writevalid_41) begin
            _saxi_register_fsm <= _saxi_register_fsm_3;
          end 
        end
        _saxi_register_fsm_1: begin
          if(saxi_rready || !saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_2;
          end 
        end
        _saxi_register_fsm_2: begin
          if(saxi_rready && saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
        _saxi_register_fsm_3: begin
          if(saxi_wvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_4;
          end 
        end
        _saxi_register_fsm_4: begin
          if(saxi_bready && saxi_bvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    _rst_logic_1 <= rst_logic;
    _rst_logic_2 <= _rst_logic_1;
    RST <= rst_logic | _rst_logic_1 | _rst_logic_2;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq <= 0;
    end else begin
      irq <= |irq_49;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_busy_edge_50 <= 0;
    end else begin
      irq_busy_edge_50 <= irq_busy;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_extern_edge_52 <= 0;
    end else begin
      irq_extern_edge_52 <= irq_extern;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_2057_1 <= 0;
      __tmp_2235_1 <= 0;
    end else begin
      __tmp_2057_1 <= _tmp_2057;
      __tmp_2235_1 <= _tmp_2235;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_2238_1 <= 0;
    end else begin
      __tmp_2238_1 <= _tmp_2238;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_2169_1 <= 0;
      __tmp_2232_1 <= 0;
    end else begin
      __tmp_2169_1 <= _tmp_2169;
      __tmp_2232_1 <= _tmp_2232;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_297_1 <= 0;
    end else begin
      __tmp_297_1 <= _tmp_297;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_300_1 <= 0;
    end else begin
      __tmp_300_1 <= _tmp_300;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_303_1 <= 0;
    end else begin
      __tmp_303_1 <= _tmp_303;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_306_1 <= 0;
    end else begin
      __tmp_306_1 <= _tmp_306;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_309_1 <= 0;
    end else begin
      __tmp_309_1 <= _tmp_309;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_312_1 <= 0;
    end else begin
      __tmp_312_1 <= _tmp_312;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_315_1 <= 0;
    end else begin
      __tmp_315_1 <= _tmp_315;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_318_1 <= 0;
    end else begin
      __tmp_318_1 <= _tmp_318;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_321_1 <= 0;
    end else begin
      __tmp_321_1 <= _tmp_321;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_2215_1 <= 0;
    end else begin
      __tmp_2215_1 <= _tmp_2215;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_2219_1 <= 0;
    end else begin
      __tmp_2219_1 <= _tmp_2219;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_324_1 <= 0;
      __tmp_2498_1 <= 0;
    end else begin
      __tmp_324_1 <= _tmp_324;
      __tmp_2498_1 <= _tmp_2498;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_327_1 <= 0;
    end else begin
      __tmp_327_1 <= _tmp_327;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_330_1 <= 0;
    end else begin
      __tmp_330_1 <= _tmp_330;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_333_1 <= 0;
    end else begin
      __tmp_333_1 <= _tmp_333;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_336_1 <= 0;
    end else begin
      __tmp_336_1 <= _tmp_336;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_339_1 <= 0;
    end else begin
      __tmp_339_1 <= _tmp_339;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_342_1 <= 0;
    end else begin
      __tmp_342_1 <= _tmp_342;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_345_1 <= 0;
    end else begin
      __tmp_345_1 <= _tmp_345;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_348_1 <= 0;
    end else begin
      __tmp_348_1 <= _tmp_348;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_351_1 <= 0;
    end else begin
      __tmp_351_1 <= _tmp_351;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_354_1 <= 0;
    end else begin
      __tmp_354_1 <= _tmp_354;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_357_1 <= 0;
    end else begin
      __tmp_357_1 <= _tmp_357;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_360_1 <= 0;
    end else begin
      __tmp_360_1 <= _tmp_360;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_363_1 <= 0;
    end else begin
      __tmp_363_1 <= _tmp_363;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_366_1 <= 0;
    end else begin
      __tmp_366_1 <= _tmp_366;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_369_1 <= 0;
    end else begin
      __tmp_369_1 <= _tmp_369;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_372_1 <= 0;
    end else begin
      __tmp_372_1 <= _tmp_372;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_375_1 <= 0;
    end else begin
      __tmp_375_1 <= _tmp_375;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_280_1 <= 0;
    end else begin
      __tmp_280_1 <= _tmp_280;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_284_1 <= 0;
    end else begin
      __tmp_284_1 <= _tmp_284;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_2043_1 <= 0;
    end else begin
      __tmp_2043_1 <= _tmp_2043;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_x_source_ram_renable <= 0;
      _acc_0_x_source_fifo_deq <= 0;
      _acc_0_x_idle <= 1;
      _acc_0_rshift_source_ram_renable <= 0;
      _acc_0_rshift_source_fifo_deq <= 0;
      _acc_0_rshift_idle <= 1;
      _acc_0_sum_sink_wenable <= 0;
      _acc_0_sum_sink_fifo_enq <= 0;
      _acc_0_valid_sink_wenable <= 0;
      _acc_0_valid_sink_fifo_enq <= 0;
      __acc_0_stream_ivalid_1 <= 0;
      __acc_0_stream_ivalid_2 <= 0;
      __acc_0_stream_ivalid_3 <= 0;
      __acc_0_stream_ivalid_4 <= 0;
      __acc_0_stream_ivalid_5 <= 0;
      _greaterthan_data_3 <= 0;
      _minus_data_5 <= 0;
      _reduceadd_data_16 <= 1'sd0;
      _reduceadd_count_16 <= 0;
      _reduceadd_prev_count_max_16 <= 0;
      _pulse_data_18 <= 1'sd0;
      _pulse_count_18 <= 0;
      _pulse_prev_count_max_18 <= 0;
      __delay_data_1964__variable_1 <= 0;
      _sll_data_7 <= 0;
      __delay_data_1961_greaterthan_3 <= 0;
      __delay_data_1962_reduceadd_16 <= 0;
      __delay_data_1965__delay_1964__variable_1 <= 0;
      __delay_data_1968_pulse_18 <= 0;
      _cond_data_13 <= 0;
      __delay_data_1963__delay_1962_reduceadd_16 <= 0;
      __delay_data_1966__delay_1965__delay_1964__variable_1 <= 0;
      __delay_data_1969__delay_1968_pulse_18 <= 0;
      _plus_data_20 <= 0;
      __delay_data_1967__delay_1966__delay_1965____variable_1 <= 0;
      __delay_data_1970__delay_1969__delay_1968_pulse_18 <= 0;
      _sra_data_21 <= 0;
      __delay_data_1971__delay_1970__delay_1969__delay_1968_pulse_18 <= 0;
      __variable_wdata_15 <= 0;
      __variable_wdata_0 <= 0;
      __variable_wdata_1 <= 0;
      __variable_wdata_2 <= 0;
      _tmp_1119 <= 0;
      _tmp_1120 <= 0;
      _tmp_1121 <= 0;
      _tmp_1122 <= 0;
      _tmp_1123 <= 0;
      _tmp_1124 <= 0;
      _tmp_1125 <= 0;
      _tmp_1126 <= 0;
      _tmp_1127 <= 0;
      _tmp_1128 <= 0;
      _tmp_1129 <= 0;
      _tmp_1130 <= 0;
      _tmp_1131 <= 0;
      _tmp_1132 <= 0;
      _tmp_1133 <= 0;
      _tmp_1134 <= 0;
      _tmp_1135 <= 0;
      _tmp_1136 <= 0;
      _tmp_1137 <= 0;
      _tmp_1138 <= 0;
      _tmp_1139 <= 0;
      _tmp_1140 <= 0;
      _tmp_1141 <= 0;
      _tmp_1142 <= 0;
      _tmp_1143 <= 0;
      _tmp_1144 <= 0;
      _tmp_1145 <= 0;
      _tmp_1146 <= 0;
      _tmp_1147 <= 0;
      _tmp_1148 <= 0;
      _tmp_1149 <= 0;
      _tmp_1150 <= 0;
      _acc_0_busy_reg <= 0;
    end else begin
      if(_acc_0_stream_oready) begin
        _acc_0_x_source_ram_renable <= 0;
        _acc_0_x_source_fifo_deq <= 0;
      end 
      _acc_0_x_idle <= _acc_0_x_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_rshift_source_ram_renable <= 0;
        _acc_0_rshift_source_fifo_deq <= 0;
      end 
      _acc_0_rshift_idle <= _acc_0_rshift_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_sum_sink_wenable <= 0;
        _acc_0_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        _acc_0_valid_sink_wenable <= 0;
        _acc_0_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_1 <= _acc_0_stream_ivalid;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_2 <= __acc_0_stream_ivalid_1;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_3 <= __acc_0_stream_ivalid_2;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_4 <= __acc_0_stream_ivalid_3;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_5 <= __acc_0_stream_ivalid_4;
      end 
      if(_acc_0_stream_oready) begin
        _greaterthan_data_3 <= acc_0_rshift_data > 1'sd0;
      end 
      if(_acc_0_stream_oready) begin
        _minus_data_5 <= acc_0_rshift_data - 2'sd1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _reduceadd_reset_cond_16) begin
        _reduceadd_data_16 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_count_16 <= (_reduceadd_current_count_16 >= acc_0_size_data - 1)? 0 : _reduceadd_current_count_16 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_prev_count_max_16 <= _reduceadd_current_count_16 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_data_16 <= _reduceadd_current_data_16 + acc_0_x_data;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _pulse_reset_cond_18) begin
        _pulse_data_18 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_count_18 <= (_pulse_current_count_18 >= acc_0_size_data - 1)? 0 : _pulse_current_count_18 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_prev_count_max_18 <= _pulse_current_count_18 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_data_18 <= _pulse_current_count_18 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1964__variable_1 <= acc_0_rshift_data;
      end 
      if(_acc_0_stream_oready) begin
        _sll_data_7 <= 2'sd1 << _minus_data_5;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1961_greaterthan_3 <= _greaterthan_data_3;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1962_reduceadd_16 <= _reduceadd_data_16;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1965__delay_1964__variable_1 <= __delay_data_1964__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1968_pulse_18 <= _pulse_data_18;
      end 
      if(_acc_0_stream_oready) begin
        _cond_data_13 <= (__delay_data_1961_greaterthan_3)? _sll_data_7 : 1'sd0;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1963__delay_1962_reduceadd_16 <= __delay_data_1962_reduceadd_16;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1966__delay_1965__delay_1964__variable_1 <= __delay_data_1965__delay_1964__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1969__delay_1968_pulse_18 <= __delay_data_1968_pulse_18;
      end 
      if(_acc_0_stream_oready) begin
        _plus_data_20 <= __delay_data_1963__delay_1962_reduceadd_16 + _cond_data_13;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1967__delay_1966__delay_1965____variable_1 <= __delay_data_1966__delay_1965__delay_1964__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1970__delay_1969__delay_1968_pulse_18 <= __delay_data_1969__delay_1968_pulse_18;
      end 
      if(_acc_0_stream_oready) begin
        _sra_data_21 <= _plus_data_20 >>> __delay_data_1967__delay_1966__delay_1965____variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_1971__delay_1970__delay_1969__delay_1968_pulse_18 <= __delay_data_1970__delay_1969__delay_1968_pulse_18;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_15 <= __delay_data_2823__delay_2822__delay_2821____variable_951;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_0 <= __substreamoutput_data_1959;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1 <= __delay_data_2838__delay_2837__delay_2836___plus_1972;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_2 <= __delay_data_2854__delay_2853__delay_2852____variable_946;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1119 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1120 <= _tmp_1119;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1121 <= _tmp_1120;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1122 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1123 <= _tmp_1122;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1124 <= _tmp_1123;
      end 
      if(_acc_0_stream_oready && _tmp_1124) begin
        __variable_wdata_15 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1125 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1126 <= _tmp_1125;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1127 <= _tmp_1126;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1128 <= _tmp_1127;
      end 
      if(_acc_0_stream_oready && _tmp_1128) begin
        __variable_wdata_15 <= 0;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        __variable_wdata_15 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1129 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1130 <= _tmp_1129;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1131 <= _tmp_1130;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1132 <= _tmp_1131;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1133 <= _tmp_1132;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1134 <= _tmp_1133;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1135 <= _tmp_1134;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1136 <= _acc_0_source_stop;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1137 <= _tmp_1136;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1138 <= _tmp_1137;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1139 <= _tmp_1138;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1140 <= _tmp_1139;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1141 <= _tmp_1140;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1142 <= _tmp_1141;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1143 <= _acc_0_source_busy;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1144 <= _tmp_1143;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1145 <= _tmp_1144;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1146 <= _tmp_1145;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1147 <= _tmp_1146;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1148 <= _tmp_1147;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1149 <= _tmp_1148;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1150 <= _acc_0_sink_busy;
      end 
      if(!_acc_0_sink_busy && _tmp_1150) begin
        _acc_0_busy_reg <= 0;
      end 
      if(_acc_0_source_busy) begin
        _acc_0_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_15 <= __delay_data_3154__delay_3153__delay_3152____variable_2450;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_0 <= __substreamoutput_data_2590;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_1 <= __delay_data_3167__delay_3166__delay_3165___plus_2592;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_2 <= __delay_data_3181__delay_3180__delay_3179____variable_2445;
      end 
    end
  end

  localparam _acc_0_fsm_1 = 1;
  localparam _acc_0_fsm_2 = 2;
  localparam _acc_0_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_fsm <= _acc_0_fsm_init;
      _acc_0_source_start <= 0;
      _acc_0_source_busy <= 0;
      _acc_0_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        _acc_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _acc_0_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_acc_0_stream_oready && _tmp_1121) begin
        _acc_0_stream_ivalid <= 1;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        _acc_0_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        _acc_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _acc_0_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_acc_0_fsm)
        _acc_0_fsm_init: begin
          if(_acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
        _acc_0_fsm_1: begin
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_source_start <= 0;
            _acc_0_source_busy <= 1;
          end 
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_2;
          end 
        end
        _acc_0_fsm_2: begin
          if(_acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_3;
          end 
        end
        _acc_0_fsm_3: begin
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_source_busy <= 0;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_fsm <= _acc_0_fsm_init;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_x_source_ram_renable <= 0;
      _acc_1_x_source_fifo_deq <= 0;
      _acc_1_x_idle <= 1;
      _acc_1_rshift_source_ram_renable <= 0;
      _acc_1_rshift_source_fifo_deq <= 0;
      _acc_1_rshift_idle <= 1;
      _acc_1_sum_sink_wenable <= 0;
      _acc_1_sum_sink_fifo_enq <= 0;
      _acc_1_valid_sink_wenable <= 0;
      _acc_1_valid_sink_fifo_enq <= 0;
      __acc_1_stream_ivalid_1 <= 0;
      __acc_1_stream_ivalid_2 <= 0;
      __acc_1_stream_ivalid_3 <= 0;
      __acc_1_stream_ivalid_4 <= 0;
      __acc_1_stream_ivalid_5 <= 0;
      _greaterthan_data_25 <= 0;
      _minus_data_27 <= 0;
      _reduceadd_data_38 <= 1'sd0;
      _reduceadd_count_38 <= 0;
      _reduceadd_prev_count_max_38 <= 0;
      _pulse_data_40 <= 1'sd0;
      _pulse_count_40 <= 0;
      _pulse_prev_count_max_40 <= 0;
      __delay_data_2382__variable_23 <= 0;
      _sll_data_29 <= 0;
      __delay_data_2379_greaterthan_25 <= 0;
      __delay_data_2380_reduceadd_38 <= 0;
      __delay_data_2383__delay_2382__variable_23 <= 0;
      __delay_data_2386_pulse_40 <= 0;
      _cond_data_35 <= 0;
      __delay_data_2381__delay_2380_reduceadd_38 <= 0;
      __delay_data_2384__delay_2383__delay_2382__variable_23 <= 0;
      __delay_data_2387__delay_2386_pulse_40 <= 0;
      _plus_data_42 <= 0;
      __delay_data_2385__delay_2384__delay_2383____variable_23 <= 0;
      __delay_data_2388__delay_2387__delay_2386_pulse_40 <= 0;
      _sra_data_43 <= 0;
      __delay_data_2389__delay_2388__delay_2387__delay_2386_pulse_40 <= 0;
      __variable_wdata_37 <= 0;
      __variable_wdata_22 <= 0;
      __variable_wdata_23 <= 0;
      __variable_wdata_24 <= 0;
      _tmp_1816 <= 0;
      _tmp_1817 <= 0;
      _tmp_1818 <= 0;
      _tmp_1819 <= 0;
      _tmp_1820 <= 0;
      _tmp_1821 <= 0;
      _tmp_1822 <= 0;
      _tmp_1823 <= 0;
      _tmp_1824 <= 0;
      _tmp_1825 <= 0;
      _tmp_1826 <= 0;
      _tmp_1827 <= 0;
      _tmp_1828 <= 0;
      _tmp_1829 <= 0;
      _tmp_1830 <= 0;
      _tmp_1831 <= 0;
      _tmp_1832 <= 0;
      _tmp_1833 <= 0;
      _tmp_1834 <= 0;
      _tmp_1835 <= 0;
      _tmp_1836 <= 0;
      _tmp_1837 <= 0;
      _tmp_1838 <= 0;
      _tmp_1839 <= 0;
      _tmp_1840 <= 0;
      _tmp_1841 <= 0;
      _tmp_1842 <= 0;
      _tmp_1843 <= 0;
      _tmp_1844 <= 0;
      _tmp_1845 <= 0;
      _tmp_1846 <= 0;
      _tmp_1847 <= 0;
      _acc_1_busy_reg <= 0;
    end else begin
      if(_acc_1_stream_oready) begin
        _acc_1_x_source_ram_renable <= 0;
        _acc_1_x_source_fifo_deq <= 0;
      end 
      _acc_1_x_idle <= _acc_1_x_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_rshift_source_ram_renable <= 0;
        _acc_1_rshift_source_fifo_deq <= 0;
      end 
      _acc_1_rshift_idle <= _acc_1_rshift_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_sum_sink_wenable <= 0;
        _acc_1_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        _acc_1_valid_sink_wenable <= 0;
        _acc_1_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_1 <= _acc_1_stream_ivalid;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_2 <= __acc_1_stream_ivalid_1;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_3 <= __acc_1_stream_ivalid_2;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_4 <= __acc_1_stream_ivalid_3;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_5 <= __acc_1_stream_ivalid_4;
      end 
      if(_acc_1_stream_oready) begin
        _greaterthan_data_25 <= acc_1_rshift_data > 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        _minus_data_27 <= acc_1_rshift_data - 2'sd1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _reduceadd_reset_cond_38) begin
        _reduceadd_data_38 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_count_38 <= (_reduceadd_current_count_38 >= acc_1_size_data - 1)? 0 : _reduceadd_current_count_38 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_prev_count_max_38 <= _reduceadd_current_count_38 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_data_38 <= _reduceadd_current_data_38 + acc_1_x_data;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _pulse_reset_cond_40) begin
        _pulse_data_40 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_count_40 <= (_pulse_current_count_40 >= acc_1_size_data - 1)? 0 : _pulse_current_count_40 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_prev_count_max_40 <= _pulse_current_count_40 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_data_40 <= _pulse_current_count_40 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2382__variable_23 <= acc_1_rshift_data;
      end 
      if(_acc_1_stream_oready) begin
        _sll_data_29 <= 2'sd1 << _minus_data_27;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2379_greaterthan_25 <= _greaterthan_data_25;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2380_reduceadd_38 <= _reduceadd_data_38;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2383__delay_2382__variable_23 <= __delay_data_2382__variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2386_pulse_40 <= _pulse_data_40;
      end 
      if(_acc_1_stream_oready) begin
        _cond_data_35 <= (__delay_data_2379_greaterthan_25)? _sll_data_29 : 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2381__delay_2380_reduceadd_38 <= __delay_data_2380_reduceadd_38;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2384__delay_2383__delay_2382__variable_23 <= __delay_data_2383__delay_2382__variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2387__delay_2386_pulse_40 <= __delay_data_2386_pulse_40;
      end 
      if(_acc_1_stream_oready) begin
        _plus_data_42 <= __delay_data_2381__delay_2380_reduceadd_38 + _cond_data_35;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2385__delay_2384__delay_2383____variable_23 <= __delay_data_2384__delay_2383__delay_2382__variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2388__delay_2387__delay_2386_pulse_40 <= __delay_data_2387__delay_2386_pulse_40;
      end 
      if(_acc_1_stream_oready) begin
        _sra_data_43 <= _plus_data_42 >>> __delay_data_2385__delay_2384__delay_2383____variable_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_2389__delay_2388__delay_2387__delay_2386_pulse_40 <= __delay_data_2388__delay_2387__delay_2386_pulse_40;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_37 <= __delay_data_2823__delay_2822__delay_2821____variable_951;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_22 <= __substreamoutput_data_2377;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_23 <= __delay_data_2959__delay_2958__delay_2957___plus_2390;
      end 
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_24 <= __delay_data_2854__delay_2853__delay_2852____variable_946;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1816 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1817 <= _tmp_1816;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1818 <= _tmp_1817;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1819 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1820 <= _tmp_1819;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1821 <= _tmp_1820;
      end 
      if(_acc_1_stream_oready && _tmp_1821) begin
        __variable_wdata_37 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1822 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1823 <= _tmp_1822;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1824 <= _tmp_1823;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1825 <= _tmp_1824;
      end 
      if(_acc_1_stream_oready && _tmp_1825) begin
        __variable_wdata_37 <= 0;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        __variable_wdata_37 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1826 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1827 <= _tmp_1826;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1828 <= _tmp_1827;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1829 <= _tmp_1828;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1830 <= _tmp_1829;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1831 <= _tmp_1830;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1832 <= _tmp_1831;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1833 <= _acc_1_source_stop;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1834 <= _tmp_1833;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1835 <= _tmp_1834;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1836 <= _tmp_1835;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1837 <= _tmp_1836;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1838 <= _tmp_1837;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1839 <= _tmp_1838;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1840 <= _acc_1_source_busy;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1841 <= _tmp_1840;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1842 <= _tmp_1841;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1843 <= _tmp_1842;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1844 <= _tmp_1843;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1845 <= _tmp_1844;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1846 <= _tmp_1845;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1847 <= _acc_1_sink_busy;
      end 
      if(!_acc_1_sink_busy && _tmp_1847) begin
        _acc_1_busy_reg <= 0;
      end 
      if(_acc_1_source_busy) begin
        _acc_1_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_37 <= __delay_data_3154__delay_3153__delay_3152____variable_2450;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_22 <= __substreamoutput_data_2621;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_23 <= __delay_data_3204__delay_3203__delay_3202___plus_2623;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_24 <= __delay_data_3181__delay_3180__delay_3179____variable_2445;
      end 
    end
  end

  localparam _acc_1_fsm_1 = 1;
  localparam _acc_1_fsm_2 = 2;
  localparam _acc_1_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_fsm <= _acc_1_fsm_init;
      _acc_1_source_start <= 0;
      _acc_1_source_busy <= 0;
      _acc_1_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_16 && _stream_conv2d_4_stream_oready) begin
        _acc_1_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _acc_1_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_acc_1_stream_oready && _tmp_1818) begin
        _acc_1_stream_ivalid <= 1;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        _acc_1_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_14 && _stream_matmul_16_stream_oready) begin
        _acc_1_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _acc_1_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_acc_1_fsm)
        _acc_1_fsm_init: begin
          if(_acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
        _acc_1_fsm_1: begin
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_source_start <= 0;
            _acc_1_source_busy <= 1;
          end 
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_2;
          end 
        end
        _acc_1_fsm_2: begin
          if(_acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_3;
          end 
        end
        _acc_1_fsm_3: begin
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_source_busy <= 0;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_fsm <= _acc_1_fsm_init;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_var0_source_ram_renable <= 0;
      _add_tree_2_var0_source_fifo_deq <= 0;
      _add_tree_2_var0_idle <= 1;
      _add_tree_2_var1_source_ram_renable <= 0;
      _add_tree_2_var1_source_fifo_deq <= 0;
      _add_tree_2_var1_idle <= 1;
      _add_tree_2_sum_sink_wenable <= 0;
      _add_tree_2_sum_sink_fifo_enq <= 0;
      __add_tree_2_stream_ivalid_1 <= 0;
      __plusn_data_47 <= 0;
      __variable_wdata_44 <= 0;
      __variable_wdata_45 <= 0;
      _tmp_2345 <= 0;
      _tmp_2346 <= 0;
      _tmp_2347 <= 0;
      _tmp_2348 <= 0;
      _tmp_2349 <= 0;
      _tmp_2350 <= 0;
      _tmp_2351 <= 0;
      _tmp_2352 <= 0;
      _tmp_2353 <= 0;
      _tmp_2354 <= 0;
      _tmp_2355 <= 0;
      _tmp_2356 <= 0;
      _tmp_2357 <= 0;
      _add_tree_2_busy_reg <= 0;
    end else begin
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var0_source_ram_renable <= 0;
        _add_tree_2_var0_source_fifo_deq <= 0;
      end 
      _add_tree_2_var0_idle <= _add_tree_2_var0_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var1_source_ram_renable <= 0;
        _add_tree_2_var1_source_fifo_deq <= 0;
      end 
      _add_tree_2_var1_idle <= _add_tree_2_var1_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_sum_sink_wenable <= 0;
        _add_tree_2_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_2_stream_oready) begin
        __add_tree_2_stream_ivalid_1 <= _add_tree_2_stream_ivalid;
      end 
      if(_add_tree_2_stream_oready) begin
        __plusn_data_47 <= add_tree_2_var0_data + add_tree_2_var1_data + 1'sd0;
      end 
      if(__stream_matmul_16_stream_ivalid_12 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_44 <= __substreamoutput_data_2583;
      end 
      if(__stream_matmul_16_stream_ivalid_12 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_45 <= __substreamoutput_data_2588;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2345 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2346 <= _tmp_2345;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2347 <= _tmp_2346;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2348 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2349 <= _tmp_2348;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2350 <= _tmp_2349;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2351 <= _add_tree_2_source_stop;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2352 <= _tmp_2351;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2353 <= _tmp_2352;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2354 <= _add_tree_2_source_busy;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2355 <= _tmp_2354;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2356 <= _tmp_2355;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_2357 <= _add_tree_2_sink_busy;
      end 
      if(!_add_tree_2_sink_busy && _tmp_2357) begin
        _add_tree_2_busy_reg <= 0;
      end 
      if(_add_tree_2_source_busy) begin
        _add_tree_2_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_2_fsm_1 = 1;
  localparam _add_tree_2_fsm_2 = 2;
  localparam _add_tree_2_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_fsm <= _add_tree_2_fsm_init;
      _add_tree_2_source_start <= 0;
      _add_tree_2_source_busy <= 0;
      _add_tree_2_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_16_stream_ivalid_12 && _stream_matmul_16_stream_oready) begin
        _add_tree_2_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _add_tree_2_source_busy <= _stream_matmul_16_source_busy;
      end 
      if(_add_tree_2_stream_oready && _tmp_2347) begin
        _add_tree_2_stream_ivalid <= 1;
      end 
      if(_add_tree_2_stream_oready && 1'd0) begin
        _add_tree_2_stream_ivalid <= 0;
      end 
      case(_add_tree_2_fsm)
        _add_tree_2_fsm_init: begin
          if(_add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
        _add_tree_2_fsm_1: begin
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_source_start <= 0;
            _add_tree_2_source_busy <= 1;
          end 
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_2;
          end 
        end
        _add_tree_2_fsm_2: begin
          if(_add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_3;
          end 
        end
        _add_tree_2_fsm_3: begin
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_source_busy <= 0;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_init;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_3_var0_source_ram_renable <= 0;
      _add_tree_3_var0_source_fifo_deq <= 0;
      _add_tree_3_var0_idle <= 1;
      _add_tree_3_var1_source_ram_renable <= 0;
      _add_tree_3_var1_source_fifo_deq <= 0;
      _add_tree_3_var1_idle <= 1;
      _add_tree_3_sum_sink_wenable <= 0;
      _add_tree_3_sum_sink_fifo_enq <= 0;
      __add_tree_3_stream_ivalid_1 <= 0;
      __plusn_data_51 <= 0;
      __variable_wdata_48 <= 0;
      __variable_wdata_49 <= 0;
      _tmp_2358 <= 0;
      _tmp_2359 <= 0;
      _tmp_2360 <= 0;
      _tmp_2361 <= 0;
      _tmp_2362 <= 0;
      _tmp_2363 <= 0;
      _tmp_2364 <= 0;
      _tmp_2365 <= 0;
      _tmp_2366 <= 0;
      _tmp_2367 <= 0;
      _tmp_2368 <= 0;
      _tmp_2369 <= 0;
      _tmp_2370 <= 0;
      _add_tree_3_busy_reg <= 0;
    end else begin
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var0_source_ram_renable <= 0;
        _add_tree_3_var0_source_fifo_deq <= 0;
      end 
      _add_tree_3_var0_idle <= _add_tree_3_var0_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var1_source_ram_renable <= 0;
        _add_tree_3_var1_source_fifo_deq <= 0;
      end 
      _add_tree_3_var1_idle <= _add_tree_3_var1_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_sum_sink_wenable <= 0;
        _add_tree_3_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_3_stream_oready) begin
        __add_tree_3_stream_ivalid_1 <= _add_tree_3_stream_ivalid;
      end 
      if(_add_tree_3_stream_oready) begin
        __plusn_data_51 <= add_tree_3_var0_data + add_tree_3_var1_data + 1'sd0;
      end 
      if(__stream_matmul_16_stream_ivalid_12 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_48 <= __substreamoutput_data_2614;
      end 
      if(__stream_matmul_16_stream_ivalid_12 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_49 <= __substreamoutput_data_2619;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2358 <= _add_tree_3_source_start;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2359 <= _tmp_2358;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2360 <= _tmp_2359;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2361 <= _add_tree_3_source_start;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2362 <= _tmp_2361;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2363 <= _tmp_2362;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2364 <= _add_tree_3_source_stop;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2365 <= _tmp_2364;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2366 <= _tmp_2365;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2367 <= _add_tree_3_source_busy;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2368 <= _tmp_2367;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2369 <= _tmp_2368;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_2370 <= _add_tree_3_sink_busy;
      end 
      if(!_add_tree_3_sink_busy && _tmp_2370) begin
        _add_tree_3_busy_reg <= 0;
      end 
      if(_add_tree_3_source_busy) begin
        _add_tree_3_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_3_fsm_1 = 1;
  localparam _add_tree_3_fsm_2 = 2;
  localparam _add_tree_3_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_3_fsm <= _add_tree_3_fsm_init;
      _add_tree_3_source_start <= 0;
      _add_tree_3_source_busy <= 0;
      _add_tree_3_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_16_stream_ivalid_12 && _stream_matmul_16_stream_oready) begin
        _add_tree_3_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _add_tree_3_source_busy <= _stream_matmul_16_source_busy;
      end 
      if(_add_tree_3_stream_oready && _tmp_2360) begin
        _add_tree_3_stream_ivalid <= 1;
      end 
      if(_add_tree_3_stream_oready && 1'd0) begin
        _add_tree_3_stream_ivalid <= 0;
      end 
      case(_add_tree_3_fsm)
        _add_tree_3_fsm_init: begin
          if(_add_tree_3_run_flag) begin
            _add_tree_3_source_start <= 1;
          end 
          if(_add_tree_3_run_flag) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_1;
          end 
        end
        _add_tree_3_fsm_1: begin
          if(_add_tree_3_source_start && _add_tree_3_stream_oready) begin
            _add_tree_3_source_start <= 0;
            _add_tree_3_source_busy <= 1;
          end 
          if(_add_tree_3_source_start && _add_tree_3_stream_oready) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_2;
          end 
        end
        _add_tree_3_fsm_2: begin
          if(_add_tree_3_stream_oready) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_3;
          end 
        end
        _add_tree_3_fsm_3: begin
          if(_add_tree_3_stream_oready && 1'd0) begin
            _add_tree_3_source_busy <= 0;
          end 
          if(_add_tree_3_stream_oready && 1'd0 && _add_tree_3_run_flag) begin
            _add_tree_3_source_start <= 1;
          end 
          if(_add_tree_3_stream_oready && 1'd0) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_init;
          end 
          if(_add_tree_3_stream_oready && 1'd0 && _add_tree_3_run_flag) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_4_var0_source_ram_renable <= 0;
      _add_tree_4_var0_source_fifo_deq <= 0;
      _add_tree_4_var0_idle <= 1;
      _add_tree_4_var1_source_ram_renable <= 0;
      _add_tree_4_var1_source_fifo_deq <= 0;
      _add_tree_4_var1_idle <= 1;
      _add_tree_4_var2_source_ram_renable <= 0;
      _add_tree_4_var2_source_fifo_deq <= 0;
      _add_tree_4_var2_idle <= 1;
      _add_tree_4_var3_source_ram_renable <= 0;
      _add_tree_4_var3_source_fifo_deq <= 0;
      _add_tree_4_var3_idle <= 1;
      _add_tree_4_var4_source_ram_renable <= 0;
      _add_tree_4_var4_source_fifo_deq <= 0;
      _add_tree_4_var4_idle <= 1;
      _add_tree_4_var5_source_ram_renable <= 0;
      _add_tree_4_var5_source_fifo_deq <= 0;
      _add_tree_4_var5_idle <= 1;
      _add_tree_4_var6_source_ram_renable <= 0;
      _add_tree_4_var6_source_fifo_deq <= 0;
      _add_tree_4_var6_idle <= 1;
      _add_tree_4_var7_source_ram_renable <= 0;
      _add_tree_4_var7_source_fifo_deq <= 0;
      _add_tree_4_var7_idle <= 1;
      _add_tree_4_var8_source_ram_renable <= 0;
      _add_tree_4_var8_source_fifo_deq <= 0;
      _add_tree_4_var8_idle <= 1;
      _add_tree_4_var9_source_ram_renable <= 0;
      _add_tree_4_var9_source_fifo_deq <= 0;
      _add_tree_4_var9_idle <= 1;
      _add_tree_4_var10_source_ram_renable <= 0;
      _add_tree_4_var10_source_fifo_deq <= 0;
      _add_tree_4_var10_idle <= 1;
      _add_tree_4_var11_source_ram_renable <= 0;
      _add_tree_4_var11_source_fifo_deq <= 0;
      _add_tree_4_var11_idle <= 1;
      _add_tree_4_var12_source_ram_renable <= 0;
      _add_tree_4_var12_source_fifo_deq <= 0;
      _add_tree_4_var12_idle <= 1;
      _add_tree_4_var13_source_ram_renable <= 0;
      _add_tree_4_var13_source_fifo_deq <= 0;
      _add_tree_4_var13_idle <= 1;
      _add_tree_4_var14_source_ram_renable <= 0;
      _add_tree_4_var14_source_fifo_deq <= 0;
      _add_tree_4_var14_idle <= 1;
      _add_tree_4_var15_source_ram_renable <= 0;
      _add_tree_4_var15_source_fifo_deq <= 0;
      _add_tree_4_var15_idle <= 1;
      _add_tree_4_var16_source_ram_renable <= 0;
      _add_tree_4_var16_source_fifo_deq <= 0;
      _add_tree_4_var16_idle <= 1;
      _add_tree_4_var17_source_ram_renable <= 0;
      _add_tree_4_var17_source_fifo_deq <= 0;
      _add_tree_4_var17_idle <= 1;
      _add_tree_4_sum_sink_wenable <= 0;
      _add_tree_4_sum_sink_fifo_enq <= 0;
      __add_tree_4_stream_ivalid_1 <= 0;
      __add_tree_4_stream_ivalid_2 <= 0;
      __add_tree_4_stream_ivalid_3 <= 0;
      __plusn_data_71 <= 0;
      __plusn_data_72 <= 0;
      __plusn_data_73 <= 0;
      __plusn_data_75 <= 0;
      __plusn_data_76 <= 0;
      __plusn_data_77 <= 0;
      __plusn_data_74 <= 0;
      __plusn_data_78 <= 0;
      __plusn_data_79 <= 0;
      __variable_wdata_52 <= 0;
      __variable_wdata_53 <= 0;
      __variable_wdata_54 <= 0;
      __variable_wdata_55 <= 0;
      __variable_wdata_56 <= 0;
      __variable_wdata_57 <= 0;
      __variable_wdata_58 <= 0;
      __variable_wdata_59 <= 0;
      __variable_wdata_60 <= 0;
      __variable_wdata_61 <= 0;
      __variable_wdata_62 <= 0;
      __variable_wdata_63 <= 0;
      __variable_wdata_64 <= 0;
      __variable_wdata_65 <= 0;
      __variable_wdata_66 <= 0;
      __variable_wdata_67 <= 0;
      __variable_wdata_68 <= 0;
      __variable_wdata_69 <= 0;
      _tmp_1100 <= 0;
      _tmp_1101 <= 0;
      _tmp_1102 <= 0;
      _tmp_1103 <= 0;
      _tmp_1104 <= 0;
      _tmp_1105 <= 0;
      _tmp_1106 <= 0;
      _tmp_1107 <= 0;
      _tmp_1108 <= 0;
      _tmp_1109 <= 0;
      _tmp_1110 <= 0;
      _tmp_1111 <= 0;
      _tmp_1112 <= 0;
      _tmp_1113 <= 0;
      _tmp_1114 <= 0;
      _tmp_1115 <= 0;
      _tmp_1116 <= 0;
      _tmp_1117 <= 0;
      _tmp_1118 <= 0;
      _add_tree_4_busy_reg <= 0;
    end else begin
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var0_source_ram_renable <= 0;
        _add_tree_4_var0_source_fifo_deq <= 0;
      end 
      _add_tree_4_var0_idle <= _add_tree_4_var0_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var1_source_ram_renable <= 0;
        _add_tree_4_var1_source_fifo_deq <= 0;
      end 
      _add_tree_4_var1_idle <= _add_tree_4_var1_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var2_source_ram_renable <= 0;
        _add_tree_4_var2_source_fifo_deq <= 0;
      end 
      _add_tree_4_var2_idle <= _add_tree_4_var2_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var3_source_ram_renable <= 0;
        _add_tree_4_var3_source_fifo_deq <= 0;
      end 
      _add_tree_4_var3_idle <= _add_tree_4_var3_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var4_source_ram_renable <= 0;
        _add_tree_4_var4_source_fifo_deq <= 0;
      end 
      _add_tree_4_var4_idle <= _add_tree_4_var4_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var5_source_ram_renable <= 0;
        _add_tree_4_var5_source_fifo_deq <= 0;
      end 
      _add_tree_4_var5_idle <= _add_tree_4_var5_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var6_source_ram_renable <= 0;
        _add_tree_4_var6_source_fifo_deq <= 0;
      end 
      _add_tree_4_var6_idle <= _add_tree_4_var6_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var7_source_ram_renable <= 0;
        _add_tree_4_var7_source_fifo_deq <= 0;
      end 
      _add_tree_4_var7_idle <= _add_tree_4_var7_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var8_source_ram_renable <= 0;
        _add_tree_4_var8_source_fifo_deq <= 0;
      end 
      _add_tree_4_var8_idle <= _add_tree_4_var8_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var9_source_ram_renable <= 0;
        _add_tree_4_var9_source_fifo_deq <= 0;
      end 
      _add_tree_4_var9_idle <= _add_tree_4_var9_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var10_source_ram_renable <= 0;
        _add_tree_4_var10_source_fifo_deq <= 0;
      end 
      _add_tree_4_var10_idle <= _add_tree_4_var10_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var11_source_ram_renable <= 0;
        _add_tree_4_var11_source_fifo_deq <= 0;
      end 
      _add_tree_4_var11_idle <= _add_tree_4_var11_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var12_source_ram_renable <= 0;
        _add_tree_4_var12_source_fifo_deq <= 0;
      end 
      _add_tree_4_var12_idle <= _add_tree_4_var12_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var13_source_ram_renable <= 0;
        _add_tree_4_var13_source_fifo_deq <= 0;
      end 
      _add_tree_4_var13_idle <= _add_tree_4_var13_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var14_source_ram_renable <= 0;
        _add_tree_4_var14_source_fifo_deq <= 0;
      end 
      _add_tree_4_var14_idle <= _add_tree_4_var14_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var15_source_ram_renable <= 0;
        _add_tree_4_var15_source_fifo_deq <= 0;
      end 
      _add_tree_4_var15_idle <= _add_tree_4_var15_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var16_source_ram_renable <= 0;
        _add_tree_4_var16_source_fifo_deq <= 0;
      end 
      _add_tree_4_var16_idle <= _add_tree_4_var16_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_var17_source_ram_renable <= 0;
        _add_tree_4_var17_source_fifo_deq <= 0;
      end 
      _add_tree_4_var17_idle <= _add_tree_4_var17_idle;
      if(_add_tree_4_stream_oready) begin
        _add_tree_4_sum_sink_wenable <= 0;
        _add_tree_4_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_4_stream_oready) begin
        __add_tree_4_stream_ivalid_1 <= _add_tree_4_stream_ivalid;
      end 
      if(_add_tree_4_stream_oready) begin
        __add_tree_4_stream_ivalid_2 <= __add_tree_4_stream_ivalid_1;
      end 
      if(_add_tree_4_stream_oready) begin
        __add_tree_4_stream_ivalid_3 <= __add_tree_4_stream_ivalid_2;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_71 <= add_tree_4_var0_data + add_tree_4_var1_data + add_tree_4_var2_data;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_72 <= add_tree_4_var3_data + add_tree_4_var4_data + add_tree_4_var5_data;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_73 <= add_tree_4_var6_data + add_tree_4_var7_data + add_tree_4_var8_data;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_75 <= add_tree_4_var9_data + add_tree_4_var10_data + add_tree_4_var11_data;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_76 <= add_tree_4_var12_data + add_tree_4_var13_data + add_tree_4_var14_data;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_77 <= add_tree_4_var15_data + add_tree_4_var16_data + add_tree_4_var17_data;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_74 <= __plusn_data_71 + __plusn_data_72 + __plusn_data_73;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_78 <= __plusn_data_75 + __plusn_data_76 + __plusn_data_77;
      end 
      if(_add_tree_4_stream_oready) begin
        __plusn_data_79 <= __plusn_data_74 + __plusn_data_78 + 1'sd0;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_52 <= __substreamoutput_data_1616;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_53 <= __substreamoutput_data_1805;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_54 <= __substreamoutput_data_1635;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_55 <= __substreamoutput_data_1824;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_56 <= __substreamoutput_data_1654;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_57 <= __substreamoutput_data_1843;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_58 <= __substreamoutput_data_1673;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_59 <= __substreamoutput_data_1862;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_60 <= __substreamoutput_data_1692;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_61 <= __substreamoutput_data_1881;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_62 <= __substreamoutput_data_1711;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_63 <= __substreamoutput_data_1900;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_64 <= __substreamoutput_data_1730;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_65 <= __substreamoutput_data_1919;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_66 <= __substreamoutput_data_1749;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_67 <= __substreamoutput_data_1938;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_68 <= __substreamoutput_data_1768;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_69 <= __substreamoutput_data_1957;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1100 <= _add_tree_4_source_start;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1101 <= _tmp_1100;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1102 <= _tmp_1101;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1103 <= _add_tree_4_source_start;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1104 <= _tmp_1103;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1105 <= _tmp_1104;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1106 <= _tmp_1105;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1107 <= _tmp_1106;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1108 <= _add_tree_4_source_stop;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1109 <= _tmp_1108;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1110 <= _tmp_1109;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1111 <= _tmp_1110;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1112 <= _tmp_1111;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1113 <= _add_tree_4_source_busy;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1114 <= _tmp_1113;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1115 <= _tmp_1114;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1116 <= _tmp_1115;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1117 <= _tmp_1116;
      end 
      if(_add_tree_4_stream_oready) begin
        _tmp_1118 <= _add_tree_4_sink_busy;
      end 
      if(!_add_tree_4_sink_busy && _tmp_1118) begin
        _add_tree_4_busy_reg <= 0;
      end 
      if(_add_tree_4_source_busy) begin
        _add_tree_4_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_4_fsm_1 = 1;
  localparam _add_tree_4_fsm_2 = 2;
  localparam _add_tree_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_4_fsm <= _add_tree_4_fsm_init;
      _add_tree_4_source_start <= 0;
      _add_tree_4_source_busy <= 0;
      _add_tree_4_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        _add_tree_4_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _add_tree_4_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_add_tree_4_stream_oready && _tmp_1102) begin
        _add_tree_4_stream_ivalid <= 1;
      end 
      if(_add_tree_4_stream_oready && 1'd0) begin
        _add_tree_4_stream_ivalid <= 0;
      end 
      case(_add_tree_4_fsm)
        _add_tree_4_fsm_init: begin
          if(_add_tree_4_run_flag) begin
            _add_tree_4_source_start <= 1;
          end 
          if(_add_tree_4_run_flag) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_1;
          end 
        end
        _add_tree_4_fsm_1: begin
          if(_add_tree_4_source_start && _add_tree_4_stream_oready) begin
            _add_tree_4_source_start <= 0;
            _add_tree_4_source_busy <= 1;
          end 
          if(_add_tree_4_source_start && _add_tree_4_stream_oready) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_2;
          end 
        end
        _add_tree_4_fsm_2: begin
          if(_add_tree_4_stream_oready) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_3;
          end 
        end
        _add_tree_4_fsm_3: begin
          if(_add_tree_4_stream_oready && 1'd0) begin
            _add_tree_4_source_busy <= 0;
          end 
          if(_add_tree_4_stream_oready && 1'd0 && _add_tree_4_run_flag) begin
            _add_tree_4_source_start <= 1;
          end 
          if(_add_tree_4_stream_oready && 1'd0) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_init;
          end 
          if(_add_tree_4_stream_oready && 1'd0 && _add_tree_4_run_flag) begin
            _add_tree_4_fsm <= _add_tree_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_5_var0_source_ram_renable <= 0;
      _add_tree_5_var0_source_fifo_deq <= 0;
      _add_tree_5_var0_idle <= 1;
      _add_tree_5_var1_source_ram_renable <= 0;
      _add_tree_5_var1_source_fifo_deq <= 0;
      _add_tree_5_var1_idle <= 1;
      _add_tree_5_var2_source_ram_renable <= 0;
      _add_tree_5_var2_source_fifo_deq <= 0;
      _add_tree_5_var2_idle <= 1;
      _add_tree_5_var3_source_ram_renable <= 0;
      _add_tree_5_var3_source_fifo_deq <= 0;
      _add_tree_5_var3_idle <= 1;
      _add_tree_5_var4_source_ram_renable <= 0;
      _add_tree_5_var4_source_fifo_deq <= 0;
      _add_tree_5_var4_idle <= 1;
      _add_tree_5_var5_source_ram_renable <= 0;
      _add_tree_5_var5_source_fifo_deq <= 0;
      _add_tree_5_var5_idle <= 1;
      _add_tree_5_var6_source_ram_renable <= 0;
      _add_tree_5_var6_source_fifo_deq <= 0;
      _add_tree_5_var6_idle <= 1;
      _add_tree_5_var7_source_ram_renable <= 0;
      _add_tree_5_var7_source_fifo_deq <= 0;
      _add_tree_5_var7_idle <= 1;
      _add_tree_5_var8_source_ram_renable <= 0;
      _add_tree_5_var8_source_fifo_deq <= 0;
      _add_tree_5_var8_idle <= 1;
      _add_tree_5_var9_source_ram_renable <= 0;
      _add_tree_5_var9_source_fifo_deq <= 0;
      _add_tree_5_var9_idle <= 1;
      _add_tree_5_var10_source_ram_renable <= 0;
      _add_tree_5_var10_source_fifo_deq <= 0;
      _add_tree_5_var10_idle <= 1;
      _add_tree_5_var11_source_ram_renable <= 0;
      _add_tree_5_var11_source_fifo_deq <= 0;
      _add_tree_5_var11_idle <= 1;
      _add_tree_5_var12_source_ram_renable <= 0;
      _add_tree_5_var12_source_fifo_deq <= 0;
      _add_tree_5_var12_idle <= 1;
      _add_tree_5_var13_source_ram_renable <= 0;
      _add_tree_5_var13_source_fifo_deq <= 0;
      _add_tree_5_var13_idle <= 1;
      _add_tree_5_var14_source_ram_renable <= 0;
      _add_tree_5_var14_source_fifo_deq <= 0;
      _add_tree_5_var14_idle <= 1;
      _add_tree_5_var15_source_ram_renable <= 0;
      _add_tree_5_var15_source_fifo_deq <= 0;
      _add_tree_5_var15_idle <= 1;
      _add_tree_5_var16_source_ram_renable <= 0;
      _add_tree_5_var16_source_fifo_deq <= 0;
      _add_tree_5_var16_idle <= 1;
      _add_tree_5_var17_source_ram_renable <= 0;
      _add_tree_5_var17_source_fifo_deq <= 0;
      _add_tree_5_var17_idle <= 1;
      _add_tree_5_sum_sink_wenable <= 0;
      _add_tree_5_sum_sink_fifo_enq <= 0;
      __add_tree_5_stream_ivalid_1 <= 0;
      __add_tree_5_stream_ivalid_2 <= 0;
      __add_tree_5_stream_ivalid_3 <= 0;
      __plusn_data_99 <= 0;
      __plusn_data_100 <= 0;
      __plusn_data_101 <= 0;
      __plusn_data_103 <= 0;
      __plusn_data_104 <= 0;
      __plusn_data_105 <= 0;
      __plusn_data_102 <= 0;
      __plusn_data_106 <= 0;
      __plusn_data_107 <= 0;
      __variable_wdata_80 <= 0;
      __variable_wdata_81 <= 0;
      __variable_wdata_82 <= 0;
      __variable_wdata_83 <= 0;
      __variable_wdata_84 <= 0;
      __variable_wdata_85 <= 0;
      __variable_wdata_86 <= 0;
      __variable_wdata_87 <= 0;
      __variable_wdata_88 <= 0;
      __variable_wdata_89 <= 0;
      __variable_wdata_90 <= 0;
      __variable_wdata_91 <= 0;
      __variable_wdata_92 <= 0;
      __variable_wdata_93 <= 0;
      __variable_wdata_94 <= 0;
      __variable_wdata_95 <= 0;
      __variable_wdata_96 <= 0;
      __variable_wdata_97 <= 0;
      _tmp_1797 <= 0;
      _tmp_1798 <= 0;
      _tmp_1799 <= 0;
      _tmp_1800 <= 0;
      _tmp_1801 <= 0;
      _tmp_1802 <= 0;
      _tmp_1803 <= 0;
      _tmp_1804 <= 0;
      _tmp_1805 <= 0;
      _tmp_1806 <= 0;
      _tmp_1807 <= 0;
      _tmp_1808 <= 0;
      _tmp_1809 <= 0;
      _tmp_1810 <= 0;
      _tmp_1811 <= 0;
      _tmp_1812 <= 0;
      _tmp_1813 <= 0;
      _tmp_1814 <= 0;
      _tmp_1815 <= 0;
      _add_tree_5_busy_reg <= 0;
    end else begin
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var0_source_ram_renable <= 0;
        _add_tree_5_var0_source_fifo_deq <= 0;
      end 
      _add_tree_5_var0_idle <= _add_tree_5_var0_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var1_source_ram_renable <= 0;
        _add_tree_5_var1_source_fifo_deq <= 0;
      end 
      _add_tree_5_var1_idle <= _add_tree_5_var1_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var2_source_ram_renable <= 0;
        _add_tree_5_var2_source_fifo_deq <= 0;
      end 
      _add_tree_5_var2_idle <= _add_tree_5_var2_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var3_source_ram_renable <= 0;
        _add_tree_5_var3_source_fifo_deq <= 0;
      end 
      _add_tree_5_var3_idle <= _add_tree_5_var3_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var4_source_ram_renable <= 0;
        _add_tree_5_var4_source_fifo_deq <= 0;
      end 
      _add_tree_5_var4_idle <= _add_tree_5_var4_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var5_source_ram_renable <= 0;
        _add_tree_5_var5_source_fifo_deq <= 0;
      end 
      _add_tree_5_var5_idle <= _add_tree_5_var5_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var6_source_ram_renable <= 0;
        _add_tree_5_var6_source_fifo_deq <= 0;
      end 
      _add_tree_5_var6_idle <= _add_tree_5_var6_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var7_source_ram_renable <= 0;
        _add_tree_5_var7_source_fifo_deq <= 0;
      end 
      _add_tree_5_var7_idle <= _add_tree_5_var7_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var8_source_ram_renable <= 0;
        _add_tree_5_var8_source_fifo_deq <= 0;
      end 
      _add_tree_5_var8_idle <= _add_tree_5_var8_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var9_source_ram_renable <= 0;
        _add_tree_5_var9_source_fifo_deq <= 0;
      end 
      _add_tree_5_var9_idle <= _add_tree_5_var9_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var10_source_ram_renable <= 0;
        _add_tree_5_var10_source_fifo_deq <= 0;
      end 
      _add_tree_5_var10_idle <= _add_tree_5_var10_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var11_source_ram_renable <= 0;
        _add_tree_5_var11_source_fifo_deq <= 0;
      end 
      _add_tree_5_var11_idle <= _add_tree_5_var11_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var12_source_ram_renable <= 0;
        _add_tree_5_var12_source_fifo_deq <= 0;
      end 
      _add_tree_5_var12_idle <= _add_tree_5_var12_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var13_source_ram_renable <= 0;
        _add_tree_5_var13_source_fifo_deq <= 0;
      end 
      _add_tree_5_var13_idle <= _add_tree_5_var13_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var14_source_ram_renable <= 0;
        _add_tree_5_var14_source_fifo_deq <= 0;
      end 
      _add_tree_5_var14_idle <= _add_tree_5_var14_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var15_source_ram_renable <= 0;
        _add_tree_5_var15_source_fifo_deq <= 0;
      end 
      _add_tree_5_var15_idle <= _add_tree_5_var15_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var16_source_ram_renable <= 0;
        _add_tree_5_var16_source_fifo_deq <= 0;
      end 
      _add_tree_5_var16_idle <= _add_tree_5_var16_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_var17_source_ram_renable <= 0;
        _add_tree_5_var17_source_fifo_deq <= 0;
      end 
      _add_tree_5_var17_idle <= _add_tree_5_var17_idle;
      if(_add_tree_5_stream_oready) begin
        _add_tree_5_sum_sink_wenable <= 0;
        _add_tree_5_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_5_stream_oready) begin
        __add_tree_5_stream_ivalid_1 <= _add_tree_5_stream_ivalid;
      end 
      if(_add_tree_5_stream_oready) begin
        __add_tree_5_stream_ivalid_2 <= __add_tree_5_stream_ivalid_1;
      end 
      if(_add_tree_5_stream_oready) begin
        __add_tree_5_stream_ivalid_3 <= __add_tree_5_stream_ivalid_2;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_99 <= add_tree_5_var0_data + add_tree_5_var1_data + add_tree_5_var2_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_100 <= add_tree_5_var3_data + add_tree_5_var4_data + add_tree_5_var5_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_101 <= add_tree_5_var6_data + add_tree_5_var7_data + add_tree_5_var8_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_103 <= add_tree_5_var9_data + add_tree_5_var10_data + add_tree_5_var11_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_104 <= add_tree_5_var12_data + add_tree_5_var13_data + add_tree_5_var14_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_105 <= add_tree_5_var15_data + add_tree_5_var16_data + add_tree_5_var17_data;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_102 <= __plusn_data_99 + __plusn_data_100 + __plusn_data_101;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_106 <= __plusn_data_103 + __plusn_data_104 + __plusn_data_105;
      end 
      if(_add_tree_5_stream_oready) begin
        __plusn_data_107 <= __plusn_data_102 + __plusn_data_106 + 1'sd0;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_80 <= __substreamoutput_data_2034;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_81 <= __substreamoutput_data_2223;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_82 <= __substreamoutput_data_2053;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_83 <= __substreamoutput_data_2242;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_84 <= __substreamoutput_data_2072;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_85 <= __substreamoutput_data_2261;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_86 <= __substreamoutput_data_2091;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_87 <= __substreamoutput_data_2280;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_88 <= __substreamoutput_data_2110;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_89 <= __substreamoutput_data_2299;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_90 <= __substreamoutput_data_2129;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_91 <= __substreamoutput_data_2318;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_92 <= __substreamoutput_data_2148;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_93 <= __substreamoutput_data_2337;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_94 <= __substreamoutput_data_2167;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_95 <= __substreamoutput_data_2356;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_96 <= __substreamoutput_data_2186;
      end 
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_97 <= __substreamoutput_data_2375;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1797 <= _add_tree_5_source_start;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1798 <= _tmp_1797;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1799 <= _tmp_1798;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1800 <= _add_tree_5_source_start;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1801 <= _tmp_1800;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1802 <= _tmp_1801;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1803 <= _tmp_1802;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1804 <= _tmp_1803;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1805 <= _add_tree_5_source_stop;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1806 <= _tmp_1805;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1807 <= _tmp_1806;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1808 <= _tmp_1807;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1809 <= _tmp_1808;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1810 <= _add_tree_5_source_busy;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1811 <= _tmp_1810;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1812 <= _tmp_1811;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1813 <= _tmp_1812;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1814 <= _tmp_1813;
      end 
      if(_add_tree_5_stream_oready) begin
        _tmp_1815 <= _add_tree_5_sink_busy;
      end 
      if(!_add_tree_5_sink_busy && _tmp_1815) begin
        _add_tree_5_busy_reg <= 0;
      end 
      if(_add_tree_5_source_busy) begin
        _add_tree_5_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_5_fsm_1 = 1;
  localparam _add_tree_5_fsm_2 = 2;
  localparam _add_tree_5_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_5_fsm <= _add_tree_5_fsm_init;
      _add_tree_5_source_start <= 0;
      _add_tree_5_source_busy <= 0;
      _add_tree_5_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_12 && _stream_conv2d_4_stream_oready) begin
        _add_tree_5_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _add_tree_5_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_add_tree_5_stream_oready && _tmp_1799) begin
        _add_tree_5_stream_ivalid <= 1;
      end 
      if(_add_tree_5_stream_oready && 1'd0) begin
        _add_tree_5_stream_ivalid <= 0;
      end 
      case(_add_tree_5_fsm)
        _add_tree_5_fsm_init: begin
          if(_add_tree_5_run_flag) begin
            _add_tree_5_source_start <= 1;
          end 
          if(_add_tree_5_run_flag) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_1;
          end 
        end
        _add_tree_5_fsm_1: begin
          if(_add_tree_5_source_start && _add_tree_5_stream_oready) begin
            _add_tree_5_source_start <= 0;
            _add_tree_5_source_busy <= 1;
          end 
          if(_add_tree_5_source_start && _add_tree_5_stream_oready) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_2;
          end 
        end
        _add_tree_5_fsm_2: begin
          if(_add_tree_5_stream_oready) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_3;
          end 
        end
        _add_tree_5_fsm_3: begin
          if(_add_tree_5_stream_oready && 1'd0) begin
            _add_tree_5_source_busy <= 0;
          end 
          if(_add_tree_5_stream_oready && 1'd0 && _add_tree_5_run_flag) begin
            _add_tree_5_source_start <= 1;
          end 
          if(_add_tree_5_stream_oready && 1'd0) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_init;
          end 
          if(_add_tree_5_stream_oready && 1'd0 && _add_tree_5_run_flag) begin
            _add_tree_5_fsm <= _add_tree_5_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_6_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_6_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_6_x_idle <= 1;
      _mul_rshift_round_clip_6_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_6_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_6_y_idle <= 1;
      _mul_rshift_round_clip_6_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_6_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_6_rshift_idle <= 1;
      _mul_rshift_round_clip_6_z_sink_wenable <= 0;
      _mul_rshift_round_clip_6_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_6_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_111 <= 0;
      __delay_data_1977_sll_117 <= 0;
      __delay_data_1981__variable_110 <= 0;
      __delay_data_1985_eq_129 <= 0;
      __delay_data_1978__delay_1977_sll_117 <= 0;
      __delay_data_1982__delay_1981__variable_110 <= 0;
      __delay_data_1986__delay_1985_eq_129 <= 0;
      __delay_data_1979__delay_1978__delay_1977_sll_117 <= 0;
      __delay_data_1983__delay_1982__delay_1981__variable_110 <= 0;
      __delay_data_1987__delay_1986__delay_1985_eq_129 <= 0;
      __delay_data_1980__delay_1979__delay_1978__delay_1977_sll_117 <= 0;
      __delay_data_1984__delay_1983__delay_1982____variable_110 <= 0;
      __delay_data_1988__delay_1987__delay_1986__delay_1985_eq_129 <= 0;
      _cond_data_130 <= 0;
      _greaterthan_data_131 <= 0;
      _lessthan_data_135 <= 0;
      _greatereq_data_139 <= 0;
      __delay_data_1989_cond_130 <= 0;
      _cond_data_133 <= 0;
      _cond_data_137 <= 0;
      __delay_data_1990_greatereq_139 <= 0;
      _cond_data_141 <= 0;
      __variable_wdata_108 <= 0;
      __variable_wdata_109 <= 0;
      __variable_wdata_110 <= 0;
      _tmp_1151 <= 0;
      _tmp_1152 <= 0;
      _tmp_1153 <= 0;
      _tmp_1154 <= 0;
      _tmp_1155 <= 0;
      _tmp_1156 <= 0;
      _tmp_1157 <= 0;
      _tmp_1158 <= 0;
      _tmp_1159 <= 0;
      _tmp_1160 <= 0;
      _tmp_1161 <= 0;
      _tmp_1162 <= 0;
      _tmp_1163 <= 0;
      _tmp_1164 <= 0;
      _tmp_1165 <= 0;
      _tmp_1166 <= 0;
      _tmp_1167 <= 0;
      _tmp_1168 <= 0;
      _tmp_1169 <= 0;
      _tmp_1170 <= 0;
      _tmp_1171 <= 0;
      _tmp_1172 <= 0;
      _tmp_1173 <= 0;
      _tmp_1174 <= 0;
      _tmp_1175 <= 0;
      _tmp_1176 <= 0;
      _tmp_1177 <= 0;
      _tmp_1178 <= 0;
      _tmp_1179 <= 0;
      _tmp_1180 <= 0;
      _tmp_1181 <= 0;
      _tmp_1182 <= 0;
      _tmp_1183 <= 0;
      _tmp_1184 <= 0;
      _mul_rshift_round_clip_6_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_6_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_6_x_idle <= _mul_rshift_round_clip_6_x_idle;
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_6_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_6_y_idle <= _mul_rshift_round_clip_6_y_idle;
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_6_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_6_rshift_idle <= _mul_rshift_round_clip_6_rshift_idle;
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _mul_rshift_round_clip_6_z_sink_wenable <= 0;
        _mul_rshift_round_clip_6_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_1 <= _mul_rshift_round_clip_6_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_2 <= __mul_rshift_round_clip_6_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_3 <= __mul_rshift_round_clip_6_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_4 <= __mul_rshift_round_clip_6_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_5 <= __mul_rshift_round_clip_6_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_6 <= __mul_rshift_round_clip_6_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_7 <= __mul_rshift_round_clip_6_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __mul_rshift_round_clip_6_stream_ivalid_8 <= __mul_rshift_round_clip_6_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _times_mul_odata_reg_111 <= _times_mul_odata_111;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1977_sll_117 <= _sll_data_117;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1981__variable_110 <= mul_rshift_round_clip_6_rshift_data;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1985_eq_129 <= _eq_data_129;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1978__delay_1977_sll_117 <= __delay_data_1977_sll_117;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1982__delay_1981__variable_110 <= __delay_data_1981__variable_110;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1986__delay_1985_eq_129 <= __delay_data_1985_eq_129;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1979__delay_1978__delay_1977_sll_117 <= __delay_data_1978__delay_1977_sll_117;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1983__delay_1982__delay_1981__variable_110 <= __delay_data_1982__delay_1981__variable_110;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1987__delay_1986__delay_1985_eq_129 <= __delay_data_1986__delay_1985_eq_129;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1980__delay_1979__delay_1978__delay_1977_sll_117 <= __delay_data_1979__delay_1978__delay_1977_sll_117;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1984__delay_1983__delay_1982____variable_110 <= __delay_data_1983__delay_1982__delay_1981__variable_110;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1988__delay_1987__delay_1986__delay_1985_eq_129 <= __delay_data_1987__delay_1986__delay_1985_eq_129;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_130 <= (__delay_data_1988__delay_1987__delay_1986__delay_1985_eq_129)? _times_data_111 : _sra_data_127;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _greaterthan_data_131 <= _cond_data_130 > 16'sd32767;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _lessthan_data_135 <= _cond_data_130 < -16'sd32767;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _greatereq_data_139 <= _cond_data_130 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1989_cond_130 <= _cond_data_130;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_133 <= (_greaterthan_data_131)? 16'sd32767 : __delay_data_1989_cond_130;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_137 <= (_lessthan_data_135)? -16'sd32767 : __delay_data_1989_cond_130;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        __delay_data_1990_greatereq_139 <= _greatereq_data_139;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _cond_data_141 <= (__delay_data_1990_greatereq_139)? _cond_data_133 : _cond_data_137;
      end 
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_108 <= _plus_data_1975;
      end 
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_109 <= __delay_data_3072__delay_3071__delay_3070__delay_3069___cond_989;
      end 
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_110 <= __delay_data_3094__delay_3093__delay_3092___plus_1991;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1151 <= _mul_rshift_round_clip_6_source_start;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1152 <= _tmp_1151;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1153 <= _tmp_1152;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1154 <= _mul_rshift_round_clip_6_source_start;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1155 <= _tmp_1154;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1156 <= _tmp_1155;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1157 <= _tmp_1156;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1158 <= _tmp_1157;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1159 <= _tmp_1158;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1160 <= _tmp_1159;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1161 <= _tmp_1160;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1162 <= _tmp_1161;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1163 <= _tmp_1162;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1164 <= _mul_rshift_round_clip_6_source_stop;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1165 <= _tmp_1164;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1166 <= _tmp_1165;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1167 <= _tmp_1166;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1168 <= _tmp_1167;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1169 <= _tmp_1168;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1170 <= _tmp_1169;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1171 <= _tmp_1170;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1172 <= _tmp_1171;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1173 <= _tmp_1172;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1174 <= _mul_rshift_round_clip_6_source_busy;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1175 <= _tmp_1174;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1176 <= _tmp_1175;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1177 <= _tmp_1176;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1178 <= _tmp_1177;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1179 <= _tmp_1178;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1180 <= _tmp_1179;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1181 <= _tmp_1180;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1182 <= _tmp_1181;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1183 <= _tmp_1182;
      end 
      if(_mul_rshift_round_clip_6_stream_oready) begin
        _tmp_1184 <= _mul_rshift_round_clip_6_sink_busy;
      end 
      if(!_mul_rshift_round_clip_6_sink_busy && _tmp_1184) begin
        _mul_rshift_round_clip_6_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_6_source_busy) begin
        _mul_rshift_round_clip_6_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_108 <= _plus_data_2595;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_109 <= __delay_data_3370__delay_3369__delay_3368___cond_2488;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_110 <= __delay_data_3390__delay_3389__delay_3388___plus_2597;
      end 
    end
  end

  localparam _mul_rshift_round_clip_6_fsm_1 = 1;
  localparam _mul_rshift_round_clip_6_fsm_2 = 2;
  localparam _mul_rshift_round_clip_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_init;
      _mul_rshift_round_clip_6_source_start <= 0;
      _mul_rshift_round_clip_6_source_busy <= 0;
      _mul_rshift_round_clip_6_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_rshift_round_clip_6_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_rshift_round_clip_6_stream_oready && _tmp_1153) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_6_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        _mul_rshift_round_clip_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _mul_rshift_round_clip_6_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_mul_rshift_round_clip_6_fsm)
        _mul_rshift_round_clip_6_fsm_init: begin
          if(_mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_1;
          end 
        end
        _mul_rshift_round_clip_6_fsm_1: begin
          if(_mul_rshift_round_clip_6_source_start && _mul_rshift_round_clip_6_stream_oready) begin
            _mul_rshift_round_clip_6_source_start <= 0;
            _mul_rshift_round_clip_6_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_6_source_start && _mul_rshift_round_clip_6_stream_oready) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_2;
          end 
        end
        _mul_rshift_round_clip_6_fsm_2: begin
          if(_mul_rshift_round_clip_6_stream_oready) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_3;
          end 
        end
        _mul_rshift_round_clip_6_fsm_3: begin
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_6_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0 && _mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_init;
          end 
          if(_mul_rshift_round_clip_6_stream_oready && 1'd0 && _mul_rshift_round_clip_6_run_flag) begin
            _mul_rshift_round_clip_6_fsm <= _mul_rshift_round_clip_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_7_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_7_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_7_x_idle <= 1;
      _mul_rshift_round_clip_7_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_7_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_7_y_idle <= 1;
      _mul_rshift_round_clip_7_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_7_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_7_rshift_idle <= 1;
      _mul_rshift_round_clip_7_z_sink_wenable <= 0;
      _mul_rshift_round_clip_7_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_7_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_145 <= 0;
      __delay_data_2395_sll_151 <= 0;
      __delay_data_2399__variable_144 <= 0;
      __delay_data_2403_eq_163 <= 0;
      __delay_data_2396__delay_2395_sll_151 <= 0;
      __delay_data_2400__delay_2399__variable_144 <= 0;
      __delay_data_2404__delay_2403_eq_163 <= 0;
      __delay_data_2397__delay_2396__delay_2395_sll_151 <= 0;
      __delay_data_2401__delay_2400__delay_2399__variable_144 <= 0;
      __delay_data_2405__delay_2404__delay_2403_eq_163 <= 0;
      __delay_data_2398__delay_2397__delay_2396__delay_2395_sll_151 <= 0;
      __delay_data_2402__delay_2401__delay_2400____variable_144 <= 0;
      __delay_data_2406__delay_2405__delay_2404__delay_2403_eq_163 <= 0;
      _cond_data_164 <= 0;
      _greaterthan_data_165 <= 0;
      _lessthan_data_169 <= 0;
      _greatereq_data_173 <= 0;
      __delay_data_2407_cond_164 <= 0;
      _cond_data_167 <= 0;
      _cond_data_171 <= 0;
      __delay_data_2408_greatereq_173 <= 0;
      _cond_data_175 <= 0;
      __variable_wdata_142 <= 0;
      __variable_wdata_143 <= 0;
      __variable_wdata_144 <= 0;
      _tmp_1848 <= 0;
      _tmp_1849 <= 0;
      _tmp_1850 <= 0;
      _tmp_1851 <= 0;
      _tmp_1852 <= 0;
      _tmp_1853 <= 0;
      _tmp_1854 <= 0;
      _tmp_1855 <= 0;
      _tmp_1856 <= 0;
      _tmp_1857 <= 0;
      _tmp_1858 <= 0;
      _tmp_1859 <= 0;
      _tmp_1860 <= 0;
      _tmp_1861 <= 0;
      _tmp_1862 <= 0;
      _tmp_1863 <= 0;
      _tmp_1864 <= 0;
      _tmp_1865 <= 0;
      _tmp_1866 <= 0;
      _tmp_1867 <= 0;
      _tmp_1868 <= 0;
      _tmp_1869 <= 0;
      _tmp_1870 <= 0;
      _tmp_1871 <= 0;
      _tmp_1872 <= 0;
      _tmp_1873 <= 0;
      _tmp_1874 <= 0;
      _tmp_1875 <= 0;
      _tmp_1876 <= 0;
      _tmp_1877 <= 0;
      _tmp_1878 <= 0;
      _tmp_1879 <= 0;
      _tmp_1880 <= 0;
      _tmp_1881 <= 0;
      _mul_rshift_round_clip_7_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_7_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_7_x_idle <= _mul_rshift_round_clip_7_x_idle;
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_7_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_7_y_idle <= _mul_rshift_round_clip_7_y_idle;
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_7_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_7_rshift_idle <= _mul_rshift_round_clip_7_rshift_idle;
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _mul_rshift_round_clip_7_z_sink_wenable <= 0;
        _mul_rshift_round_clip_7_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_1 <= _mul_rshift_round_clip_7_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_2 <= __mul_rshift_round_clip_7_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_3 <= __mul_rshift_round_clip_7_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_4 <= __mul_rshift_round_clip_7_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_5 <= __mul_rshift_round_clip_7_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_6 <= __mul_rshift_round_clip_7_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_7 <= __mul_rshift_round_clip_7_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __mul_rshift_round_clip_7_stream_ivalid_8 <= __mul_rshift_round_clip_7_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _times_mul_odata_reg_145 <= _times_mul_odata_145;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2395_sll_151 <= _sll_data_151;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2399__variable_144 <= mul_rshift_round_clip_7_rshift_data;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2403_eq_163 <= _eq_data_163;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2396__delay_2395_sll_151 <= __delay_data_2395_sll_151;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2400__delay_2399__variable_144 <= __delay_data_2399__variable_144;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2404__delay_2403_eq_163 <= __delay_data_2403_eq_163;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2397__delay_2396__delay_2395_sll_151 <= __delay_data_2396__delay_2395_sll_151;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2401__delay_2400__delay_2399__variable_144 <= __delay_data_2400__delay_2399__variable_144;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2405__delay_2404__delay_2403_eq_163 <= __delay_data_2404__delay_2403_eq_163;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2398__delay_2397__delay_2396__delay_2395_sll_151 <= __delay_data_2397__delay_2396__delay_2395_sll_151;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2402__delay_2401__delay_2400____variable_144 <= __delay_data_2401__delay_2400__delay_2399__variable_144;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2406__delay_2405__delay_2404__delay_2403_eq_163 <= __delay_data_2405__delay_2404__delay_2403_eq_163;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_164 <= (__delay_data_2406__delay_2405__delay_2404__delay_2403_eq_163)? _times_data_145 : _sra_data_161;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _greaterthan_data_165 <= _cond_data_164 > 16'sd32767;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _lessthan_data_169 <= _cond_data_164 < -16'sd32767;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _greatereq_data_173 <= _cond_data_164 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2407_cond_164 <= _cond_data_164;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_167 <= (_greaterthan_data_165)? 16'sd32767 : __delay_data_2407_cond_164;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_171 <= (_lessthan_data_169)? -16'sd32767 : __delay_data_2407_cond_164;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        __delay_data_2408_greatereq_173 <= _greatereq_data_173;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _cond_data_175 <= (__delay_data_2408_greatereq_173)? _cond_data_167 : _cond_data_171;
      end 
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_142 <= _plus_data_2393;
      end 
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_143 <= __delay_data_3004__delay_3003__delay_3002__delay_3001___cond_990;
      end 
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_144 <= __delay_data_3026__delay_3025__delay_3024___plus_2409;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1848 <= _mul_rshift_round_clip_7_source_start;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1849 <= _tmp_1848;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1850 <= _tmp_1849;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1851 <= _mul_rshift_round_clip_7_source_start;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1852 <= _tmp_1851;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1853 <= _tmp_1852;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1854 <= _tmp_1853;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1855 <= _tmp_1854;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1856 <= _tmp_1855;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1857 <= _tmp_1856;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1858 <= _tmp_1857;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1859 <= _tmp_1858;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1860 <= _tmp_1859;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1861 <= _mul_rshift_round_clip_7_source_stop;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1862 <= _tmp_1861;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1863 <= _tmp_1862;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1864 <= _tmp_1863;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1865 <= _tmp_1864;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1866 <= _tmp_1865;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1867 <= _tmp_1866;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1868 <= _tmp_1867;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1869 <= _tmp_1868;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1870 <= _tmp_1869;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1871 <= _mul_rshift_round_clip_7_source_busy;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1872 <= _tmp_1871;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1873 <= _tmp_1872;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1874 <= _tmp_1873;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1875 <= _tmp_1874;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1876 <= _tmp_1875;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1877 <= _tmp_1876;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1878 <= _tmp_1877;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1879 <= _tmp_1878;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1880 <= _tmp_1879;
      end 
      if(_mul_rshift_round_clip_7_stream_oready) begin
        _tmp_1881 <= _mul_rshift_round_clip_7_sink_busy;
      end 
      if(!_mul_rshift_round_clip_7_sink_busy && _tmp_1881) begin
        _mul_rshift_round_clip_7_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_7_source_busy) begin
        _mul_rshift_round_clip_7_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_142 <= _plus_data_2626;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_143 <= __delay_data_3245__delay_3244__delay_3243___cond_2489;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_144 <= __delay_data_3265__delay_3264__delay_3263___plus_2628;
      end 
    end
  end

  localparam _mul_rshift_round_clip_7_fsm_1 = 1;
  localparam _mul_rshift_round_clip_7_fsm_2 = 2;
  localparam _mul_rshift_round_clip_7_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_init;
      _mul_rshift_round_clip_7_source_start <= 0;
      _mul_rshift_round_clip_7_source_busy <= 0;
      _mul_rshift_round_clip_7_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_23 && _stream_conv2d_4_stream_oready) begin
        _mul_rshift_round_clip_7_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_rshift_round_clip_7_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_rshift_round_clip_7_stream_oready && _tmp_1850) begin
        _mul_rshift_round_clip_7_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_7_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_7_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_21 && _stream_matmul_16_stream_oready) begin
        _mul_rshift_round_clip_7_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _mul_rshift_round_clip_7_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_mul_rshift_round_clip_7_fsm)
        _mul_rshift_round_clip_7_fsm_init: begin
          if(_mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_1;
          end 
        end
        _mul_rshift_round_clip_7_fsm_1: begin
          if(_mul_rshift_round_clip_7_source_start && _mul_rshift_round_clip_7_stream_oready) begin
            _mul_rshift_round_clip_7_source_start <= 0;
            _mul_rshift_round_clip_7_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_7_source_start && _mul_rshift_round_clip_7_stream_oready) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_2;
          end 
        end
        _mul_rshift_round_clip_7_fsm_2: begin
          if(_mul_rshift_round_clip_7_stream_oready) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_3;
          end 
        end
        _mul_rshift_round_clip_7_fsm_3: begin
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_7_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0 && _mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_init;
          end 
          if(_mul_rshift_round_clip_7_stream_oready && 1'd0 && _mul_rshift_round_clip_7_run_flag) begin
            _mul_rshift_round_clip_7_fsm <= _mul_rshift_round_clip_7_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_x_source_ram_renable <= 0;
      _mul_8_x_source_fifo_deq <= 0;
      _mul_8_x_idle <= 1;
      _mul_8_y_source_ram_renable <= 0;
      _mul_8_y_source_fifo_deq <= 0;
      _mul_8_y_idle <= 1;
      _mul_8_rshift_source_ram_renable <= 0;
      _mul_8_rshift_source_fifo_deq <= 0;
      _mul_8_rshift_idle <= 1;
      _mul_8_z_sink_wenable <= 0;
      _mul_8_z_sink_fifo_enq <= 0;
      __mul_8_stream_ivalid_1 <= 0;
      __mul_8_stream_ivalid_2 <= 0;
      __mul_8_stream_ivalid_3 <= 0;
      __mul_8_stream_ivalid_4 <= 0;
      __mul_8_stream_ivalid_5 <= 0;
      __mul_8_stream_ivalid_6 <= 0;
      __mul_8_stream_ivalid_7 <= 0;
      __mul_8_stream_ivalid_8 <= 0;
      _greaterthan_data_179 <= 0;
      _minus_data_181 <= 0;
      _greatereq_data_192 <= 0;
      __delay_data_1602__variable_176 <= 0;
      __delay_data_1605__variable_177 <= 0;
      __delay_data_1608__variable_178 <= 0;
      _sll_data_183 <= 0;
      __delay_data_1599_greaterthan_179 <= 0;
      __delay_data_1600_greatereq_192 <= 0;
      __delay_data_1603__delay_1602__variable_176 <= 0;
      __delay_data_1606__delay_1605__variable_177 <= 0;
      __delay_data_1609__delay_1608__variable_178 <= 0;
      _cond_data_189 <= 0;
      __delay_data_1601__delay_1600_greatereq_192 <= 0;
      __delay_data_1604__delay_1603__delay_1602__variable_176 <= 0;
      __delay_data_1607__delay_1606__delay_1605__variable_177 <= 0;
      __delay_data_1610__delay_1609__delay_1608__variable_178 <= 0;
      __muladd_madd_odata_reg_195 <= 0;
      __delay_data_1611__delay_1610__delay_1609____variable_178 <= 0;
      __delay_data_1612__delay_1611__delay_1610____variable_178 <= 0;
      __delay_data_1613__delay_1612__delay_1611____variable_178 <= 0;
      __delay_data_1614__delay_1613__delay_1612____variable_178 <= 0;
      _sra_data_196 <= 0;
      __variable_wdata_176 <= 0;
      __variable_wdata_177 <= 0;
      __variable_wdata_178 <= 0;
      _tmp_488 <= 0;
      _tmp_489 <= 0;
      _tmp_490 <= 0;
      _tmp_491 <= 0;
      _tmp_492 <= 0;
      _tmp_493 <= 0;
      _tmp_494 <= 0;
      _tmp_495 <= 0;
      _tmp_496 <= 0;
      _tmp_497 <= 0;
      _tmp_498 <= 0;
      _tmp_499 <= 0;
      _tmp_500 <= 0;
      _tmp_501 <= 0;
      _tmp_502 <= 0;
      _tmp_503 <= 0;
      _tmp_504 <= 0;
      _tmp_505 <= 0;
      _tmp_506 <= 0;
      _tmp_507 <= 0;
      _tmp_508 <= 0;
      _tmp_509 <= 0;
      _tmp_510 <= 0;
      _tmp_511 <= 0;
      _tmp_512 <= 0;
      _tmp_513 <= 0;
      _tmp_514 <= 0;
      _tmp_515 <= 0;
      _tmp_516 <= 0;
      _tmp_517 <= 0;
      _tmp_518 <= 0;
      _tmp_519 <= 0;
      _tmp_520 <= 0;
      _tmp_521 <= 0;
      _mul_8_busy_reg <= 0;
    end else begin
      if(_mul_8_stream_oready) begin
        _mul_8_x_source_ram_renable <= 0;
        _mul_8_x_source_fifo_deq <= 0;
      end 
      _mul_8_x_idle <= _mul_8_x_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_y_source_ram_renable <= 0;
        _mul_8_y_source_fifo_deq <= 0;
      end 
      _mul_8_y_idle <= _mul_8_y_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_rshift_source_ram_renable <= 0;
        _mul_8_rshift_source_fifo_deq <= 0;
      end 
      _mul_8_rshift_idle <= _mul_8_rshift_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_z_sink_wenable <= 0;
        _mul_8_z_sink_fifo_enq <= 0;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_1 <= _mul_8_stream_ivalid;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_2 <= __mul_8_stream_ivalid_1;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_3 <= __mul_8_stream_ivalid_2;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_4 <= __mul_8_stream_ivalid_3;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_5 <= __mul_8_stream_ivalid_4;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_6 <= __mul_8_stream_ivalid_5;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_7 <= __mul_8_stream_ivalid_6;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_8 <= __mul_8_stream_ivalid_7;
      end 
      if(_mul_8_stream_oready) begin
        _greaterthan_data_179 <= mul_8_rshift_data > 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        _minus_data_181 <= mul_8_rshift_data - 2'sd1;
      end 
      if(_mul_8_stream_oready) begin
        _greatereq_data_192 <= mul_8_x_data >= 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1602__variable_176 <= mul_8_x_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1605__variable_177 <= mul_8_y_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1608__variable_178 <= mul_8_rshift_data;
      end 
      if(_mul_8_stream_oready) begin
        _sll_data_183 <= 2'sd1 << _minus_data_181;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1599_greaterthan_179 <= _greaterthan_data_179;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1600_greatereq_192 <= _greatereq_data_192;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1603__delay_1602__variable_176 <= __delay_data_1602__variable_176;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1606__delay_1605__variable_177 <= __delay_data_1605__variable_177;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1609__delay_1608__variable_178 <= __delay_data_1608__variable_178;
      end 
      if(_mul_8_stream_oready) begin
        _cond_data_189 <= (__delay_data_1599_greaterthan_179)? _sll_data_183 : 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1601__delay_1600_greatereq_192 <= __delay_data_1600_greatereq_192;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1604__delay_1603__delay_1602__variable_176 <= __delay_data_1603__delay_1602__variable_176;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1607__delay_1606__delay_1605__variable_177 <= __delay_data_1606__delay_1605__variable_177;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1610__delay_1609__delay_1608__variable_178 <= __delay_data_1609__delay_1608__variable_178;
      end 
      if(_mul_8_stream_oready) begin
        __muladd_madd_odata_reg_195 <= __muladd_madd_odata_195;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1611__delay_1610__delay_1609____variable_178 <= __delay_data_1610__delay_1609__delay_1608__variable_178;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1612__delay_1611__delay_1610____variable_178 <= __delay_data_1611__delay_1610__delay_1609____variable_178;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1613__delay_1612__delay_1611____variable_178 <= __delay_data_1612__delay_1611__delay_1610____variable_178;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_1614__delay_1613__delay_1612____variable_178 <= __delay_data_1613__delay_1612__delay_1611____variable_178;
      end 
      if(_mul_8_stream_oready) begin
        _sra_data_196 <= __muladd_data_195 >>> __delay_data_1614__delay_1613__delay_1612____variable_178;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_176 <= _cond_data_1581;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_177 <= _cond_data_1419;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_178 <= __delay_data_2662__delay_2661_plus_1615;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_488 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_489 <= _tmp_488;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_490 <= _tmp_489;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_491 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_492 <= _tmp_491;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_493 <= _tmp_492;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_494 <= _tmp_493;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_495 <= _tmp_494;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_496 <= _tmp_495;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_497 <= _tmp_496;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_498 <= _tmp_497;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_499 <= _tmp_498;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_500 <= _tmp_499;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_501 <= _mul_8_source_stop;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_502 <= _tmp_501;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_503 <= _tmp_502;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_504 <= _tmp_503;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_505 <= _tmp_504;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_506 <= _tmp_505;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_507 <= _tmp_506;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_508 <= _tmp_507;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_509 <= _tmp_508;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_510 <= _tmp_509;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_511 <= _mul_8_source_busy;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_512 <= _tmp_511;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_513 <= _tmp_512;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_514 <= _tmp_513;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_515 <= _tmp_514;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_516 <= _tmp_515;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_517 <= _tmp_516;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_518 <= _tmp_517;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_519 <= _tmp_518;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_520 <= _tmp_519;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_521 <= _mul_8_sink_busy;
      end 
      if(!_mul_8_sink_busy && _tmp_521) begin
        _mul_8_busy_reg <= 0;
      end 
      if(_mul_8_source_busy) begin
        _mul_8_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_176 <= _cond_data_2580;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_177 <= _cond_data_2562;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_178 <= __delay_data_3131__delay_3130_plus_2582;
      end 
    end
  end

  localparam _mul_8_fsm_1 = 1;
  localparam _mul_8_fsm_2 = 2;
  localparam _mul_8_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_fsm <= _mul_8_fsm_init;
      _mul_8_source_start <= 0;
      _mul_8_source_busy <= 0;
      _mul_8_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_8_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_8_stream_oready && _tmp_490) begin
        _mul_8_stream_ivalid <= 1;
      end 
      if(_mul_8_stream_oready && 1'd0) begin
        _mul_8_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _mul_8_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_mul_8_fsm)
        _mul_8_fsm_init: begin
          if(_mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
        _mul_8_fsm_1: begin
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_source_start <= 0;
            _mul_8_source_busy <= 1;
          end 
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_2;
          end 
        end
        _mul_8_fsm_2: begin
          if(_mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_3;
          end 
        end
        _mul_8_fsm_3: begin
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_source_busy <= 0;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_fsm <= _mul_8_fsm_init;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_x_source_ram_renable <= 0;
      _mul_9_x_source_fifo_deq <= 0;
      _mul_9_x_idle <= 1;
      _mul_9_y_source_ram_renable <= 0;
      _mul_9_y_source_fifo_deq <= 0;
      _mul_9_y_idle <= 1;
      _mul_9_rshift_source_ram_renable <= 0;
      _mul_9_rshift_source_fifo_deq <= 0;
      _mul_9_rshift_idle <= 1;
      _mul_9_z_sink_wenable <= 0;
      _mul_9_z_sink_fifo_enq <= 0;
      __mul_9_stream_ivalid_1 <= 0;
      __mul_9_stream_ivalid_2 <= 0;
      __mul_9_stream_ivalid_3 <= 0;
      __mul_9_stream_ivalid_4 <= 0;
      __mul_9_stream_ivalid_5 <= 0;
      __mul_9_stream_ivalid_6 <= 0;
      __mul_9_stream_ivalid_7 <= 0;
      __mul_9_stream_ivalid_8 <= 0;
      _greaterthan_data_200 <= 0;
      _minus_data_202 <= 0;
      _greatereq_data_213 <= 0;
      __delay_data_1621__variable_197 <= 0;
      __delay_data_1624__variable_198 <= 0;
      __delay_data_1627__variable_199 <= 0;
      _sll_data_204 <= 0;
      __delay_data_1618_greaterthan_200 <= 0;
      __delay_data_1619_greatereq_213 <= 0;
      __delay_data_1622__delay_1621__variable_197 <= 0;
      __delay_data_1625__delay_1624__variable_198 <= 0;
      __delay_data_1628__delay_1627__variable_199 <= 0;
      _cond_data_210 <= 0;
      __delay_data_1620__delay_1619_greatereq_213 <= 0;
      __delay_data_1623__delay_1622__delay_1621__variable_197 <= 0;
      __delay_data_1626__delay_1625__delay_1624__variable_198 <= 0;
      __delay_data_1629__delay_1628__delay_1627__variable_199 <= 0;
      __muladd_madd_odata_reg_216 <= 0;
      __delay_data_1630__delay_1629__delay_1628____variable_199 <= 0;
      __delay_data_1631__delay_1630__delay_1629____variable_199 <= 0;
      __delay_data_1632__delay_1631__delay_1630____variable_199 <= 0;
      __delay_data_1633__delay_1632__delay_1631____variable_199 <= 0;
      _sra_data_217 <= 0;
      __variable_wdata_197 <= 0;
      __variable_wdata_198 <= 0;
      __variable_wdata_199 <= 0;
      _tmp_522 <= 0;
      _tmp_523 <= 0;
      _tmp_524 <= 0;
      _tmp_525 <= 0;
      _tmp_526 <= 0;
      _tmp_527 <= 0;
      _tmp_528 <= 0;
      _tmp_529 <= 0;
      _tmp_530 <= 0;
      _tmp_531 <= 0;
      _tmp_532 <= 0;
      _tmp_533 <= 0;
      _tmp_534 <= 0;
      _tmp_535 <= 0;
      _tmp_536 <= 0;
      _tmp_537 <= 0;
      _tmp_538 <= 0;
      _tmp_539 <= 0;
      _tmp_540 <= 0;
      _tmp_541 <= 0;
      _tmp_542 <= 0;
      _tmp_543 <= 0;
      _tmp_544 <= 0;
      _tmp_545 <= 0;
      _tmp_546 <= 0;
      _tmp_547 <= 0;
      _tmp_548 <= 0;
      _tmp_549 <= 0;
      _tmp_550 <= 0;
      _tmp_551 <= 0;
      _tmp_552 <= 0;
      _tmp_553 <= 0;
      _tmp_554 <= 0;
      _tmp_555 <= 0;
      _mul_9_busy_reg <= 0;
    end else begin
      if(_mul_9_stream_oready) begin
        _mul_9_x_source_ram_renable <= 0;
        _mul_9_x_source_fifo_deq <= 0;
      end 
      _mul_9_x_idle <= _mul_9_x_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_y_source_ram_renable <= 0;
        _mul_9_y_source_fifo_deq <= 0;
      end 
      _mul_9_y_idle <= _mul_9_y_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_rshift_source_ram_renable <= 0;
        _mul_9_rshift_source_fifo_deq <= 0;
      end 
      _mul_9_rshift_idle <= _mul_9_rshift_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_z_sink_wenable <= 0;
        _mul_9_z_sink_fifo_enq <= 0;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_1 <= _mul_9_stream_ivalid;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_2 <= __mul_9_stream_ivalid_1;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_3 <= __mul_9_stream_ivalid_2;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_4 <= __mul_9_stream_ivalid_3;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_5 <= __mul_9_stream_ivalid_4;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_6 <= __mul_9_stream_ivalid_5;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_7 <= __mul_9_stream_ivalid_6;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_8 <= __mul_9_stream_ivalid_7;
      end 
      if(_mul_9_stream_oready) begin
        _greaterthan_data_200 <= mul_9_rshift_data > 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        _minus_data_202 <= mul_9_rshift_data - 2'sd1;
      end 
      if(_mul_9_stream_oready) begin
        _greatereq_data_213 <= mul_9_x_data >= 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1621__variable_197 <= mul_9_x_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1624__variable_198 <= mul_9_y_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1627__variable_199 <= mul_9_rshift_data;
      end 
      if(_mul_9_stream_oready) begin
        _sll_data_204 <= 2'sd1 << _minus_data_202;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1618_greaterthan_200 <= _greaterthan_data_200;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1619_greatereq_213 <= _greatereq_data_213;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1622__delay_1621__variable_197 <= __delay_data_1621__variable_197;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1625__delay_1624__variable_198 <= __delay_data_1624__variable_198;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1628__delay_1627__variable_199 <= __delay_data_1627__variable_199;
      end 
      if(_mul_9_stream_oready) begin
        _cond_data_210 <= (__delay_data_1618_greaterthan_200)? _sll_data_204 : 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1620__delay_1619_greatereq_213 <= __delay_data_1619_greatereq_213;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1623__delay_1622__delay_1621__variable_197 <= __delay_data_1622__delay_1621__variable_197;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1626__delay_1625__delay_1624__variable_198 <= __delay_data_1625__delay_1624__variable_198;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1629__delay_1628__delay_1627__variable_199 <= __delay_data_1628__delay_1627__variable_199;
      end 
      if(_mul_9_stream_oready) begin
        __muladd_madd_odata_reg_216 <= __muladd_madd_odata_216;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1630__delay_1629__delay_1628____variable_199 <= __delay_data_1629__delay_1628__delay_1627__variable_199;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1631__delay_1630__delay_1629____variable_199 <= __delay_data_1630__delay_1629__delay_1628____variable_199;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1632__delay_1631__delay_1630____variable_199 <= __delay_data_1631__delay_1630__delay_1629____variable_199;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_1633__delay_1632__delay_1631____variable_199 <= __delay_data_1632__delay_1631__delay_1630____variable_199;
      end 
      if(_mul_9_stream_oready) begin
        _sra_data_217 <= __muladd_data_216 >>> __delay_data_1633__delay_1632__delay_1631____variable_199;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_197 <= _cond_data_1583;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_198 <= _cond_data_1421;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_199 <= __delay_data_2681__delay_2680_plus_1634;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_522 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_523 <= _tmp_522;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_524 <= _tmp_523;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_525 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_526 <= _tmp_525;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_527 <= _tmp_526;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_528 <= _tmp_527;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_529 <= _tmp_528;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_530 <= _tmp_529;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_531 <= _tmp_530;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_532 <= _tmp_531;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_533 <= _tmp_532;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_534 <= _tmp_533;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_535 <= _mul_9_source_stop;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_536 <= _tmp_535;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_537 <= _tmp_536;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_538 <= _tmp_537;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_539 <= _tmp_538;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_540 <= _tmp_539;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_541 <= _tmp_540;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_542 <= _tmp_541;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_543 <= _tmp_542;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_544 <= _tmp_543;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_545 <= _mul_9_source_busy;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_546 <= _tmp_545;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_547 <= _tmp_546;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_548 <= _tmp_547;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_549 <= _tmp_548;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_550 <= _tmp_549;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_551 <= _tmp_550;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_552 <= _tmp_551;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_553 <= _tmp_552;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_554 <= _tmp_553;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_555 <= _mul_9_sink_busy;
      end 
      if(!_mul_9_sink_busy && _tmp_555) begin
        _mul_9_busy_reg <= 0;
      end 
      if(_mul_9_source_busy) begin
        _mul_9_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_197 <= _cond_data_2585;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_198 <= _cond_data_2564;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_199 <= __delay_data_3140__delay_3139_plus_2587;
      end 
    end
  end

  localparam _mul_9_fsm_1 = 1;
  localparam _mul_9_fsm_2 = 2;
  localparam _mul_9_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_fsm <= _mul_9_fsm_init;
      _mul_9_source_start <= 0;
      _mul_9_source_busy <= 0;
      _mul_9_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_9_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_9_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_9_stream_oready && _tmp_524) begin
        _mul_9_stream_ivalid <= 1;
      end 
      if(_mul_9_stream_oready && 1'd0) begin
        _mul_9_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        _mul_9_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _mul_9_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_mul_9_fsm)
        _mul_9_fsm_init: begin
          if(_mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
        _mul_9_fsm_1: begin
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_source_start <= 0;
            _mul_9_source_busy <= 1;
          end 
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_2;
          end 
        end
        _mul_9_fsm_2: begin
          if(_mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_3;
          end 
        end
        _mul_9_fsm_3: begin
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_source_busy <= 0;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_fsm <= _mul_9_fsm_init;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_x_source_ram_renable <= 0;
      _mul_10_x_source_fifo_deq <= 0;
      _mul_10_x_idle <= 1;
      _mul_10_y_source_ram_renable <= 0;
      _mul_10_y_source_fifo_deq <= 0;
      _mul_10_y_idle <= 1;
      _mul_10_rshift_source_ram_renable <= 0;
      _mul_10_rshift_source_fifo_deq <= 0;
      _mul_10_rshift_idle <= 1;
      _mul_10_z_sink_wenable <= 0;
      _mul_10_z_sink_fifo_enq <= 0;
      __mul_10_stream_ivalid_1 <= 0;
      __mul_10_stream_ivalid_2 <= 0;
      __mul_10_stream_ivalid_3 <= 0;
      __mul_10_stream_ivalid_4 <= 0;
      __mul_10_stream_ivalid_5 <= 0;
      __mul_10_stream_ivalid_6 <= 0;
      __mul_10_stream_ivalid_7 <= 0;
      __mul_10_stream_ivalid_8 <= 0;
      _greaterthan_data_221 <= 0;
      _minus_data_223 <= 0;
      _greatereq_data_234 <= 0;
      __delay_data_1640__variable_218 <= 0;
      __delay_data_1643__variable_219 <= 0;
      __delay_data_1646__variable_220 <= 0;
      _sll_data_225 <= 0;
      __delay_data_1637_greaterthan_221 <= 0;
      __delay_data_1638_greatereq_234 <= 0;
      __delay_data_1641__delay_1640__variable_218 <= 0;
      __delay_data_1644__delay_1643__variable_219 <= 0;
      __delay_data_1647__delay_1646__variable_220 <= 0;
      _cond_data_231 <= 0;
      __delay_data_1639__delay_1638_greatereq_234 <= 0;
      __delay_data_1642__delay_1641__delay_1640__variable_218 <= 0;
      __delay_data_1645__delay_1644__delay_1643__variable_219 <= 0;
      __delay_data_1648__delay_1647__delay_1646__variable_220 <= 0;
      __muladd_madd_odata_reg_237 <= 0;
      __delay_data_1649__delay_1648__delay_1647____variable_220 <= 0;
      __delay_data_1650__delay_1649__delay_1648____variable_220 <= 0;
      __delay_data_1651__delay_1650__delay_1649____variable_220 <= 0;
      __delay_data_1652__delay_1651__delay_1650____variable_220 <= 0;
      _sra_data_238 <= 0;
      __variable_wdata_218 <= 0;
      __variable_wdata_219 <= 0;
      __variable_wdata_220 <= 0;
      _tmp_556 <= 0;
      _tmp_557 <= 0;
      _tmp_558 <= 0;
      _tmp_559 <= 0;
      _tmp_560 <= 0;
      _tmp_561 <= 0;
      _tmp_562 <= 0;
      _tmp_563 <= 0;
      _tmp_564 <= 0;
      _tmp_565 <= 0;
      _tmp_566 <= 0;
      _tmp_567 <= 0;
      _tmp_568 <= 0;
      _tmp_569 <= 0;
      _tmp_570 <= 0;
      _tmp_571 <= 0;
      _tmp_572 <= 0;
      _tmp_573 <= 0;
      _tmp_574 <= 0;
      _tmp_575 <= 0;
      _tmp_576 <= 0;
      _tmp_577 <= 0;
      _tmp_578 <= 0;
      _tmp_579 <= 0;
      _tmp_580 <= 0;
      _tmp_581 <= 0;
      _tmp_582 <= 0;
      _tmp_583 <= 0;
      _tmp_584 <= 0;
      _tmp_585 <= 0;
      _tmp_586 <= 0;
      _tmp_587 <= 0;
      _tmp_588 <= 0;
      _tmp_589 <= 0;
      _mul_10_busy_reg <= 0;
    end else begin
      if(_mul_10_stream_oready) begin
        _mul_10_x_source_ram_renable <= 0;
        _mul_10_x_source_fifo_deq <= 0;
      end 
      _mul_10_x_idle <= _mul_10_x_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_y_source_ram_renable <= 0;
        _mul_10_y_source_fifo_deq <= 0;
      end 
      _mul_10_y_idle <= _mul_10_y_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_rshift_source_ram_renable <= 0;
        _mul_10_rshift_source_fifo_deq <= 0;
      end 
      _mul_10_rshift_idle <= _mul_10_rshift_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_z_sink_wenable <= 0;
        _mul_10_z_sink_fifo_enq <= 0;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_1 <= _mul_10_stream_ivalid;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_2 <= __mul_10_stream_ivalid_1;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_3 <= __mul_10_stream_ivalid_2;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_4 <= __mul_10_stream_ivalid_3;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_5 <= __mul_10_stream_ivalid_4;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_6 <= __mul_10_stream_ivalid_5;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_7 <= __mul_10_stream_ivalid_6;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_8 <= __mul_10_stream_ivalid_7;
      end 
      if(_mul_10_stream_oready) begin
        _greaterthan_data_221 <= mul_10_rshift_data > 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        _minus_data_223 <= mul_10_rshift_data - 2'sd1;
      end 
      if(_mul_10_stream_oready) begin
        _greatereq_data_234 <= mul_10_x_data >= 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1640__variable_218 <= mul_10_x_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1643__variable_219 <= mul_10_y_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1646__variable_220 <= mul_10_rshift_data;
      end 
      if(_mul_10_stream_oready) begin
        _sll_data_225 <= 2'sd1 << _minus_data_223;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1637_greaterthan_221 <= _greaterthan_data_221;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1638_greatereq_234 <= _greatereq_data_234;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1641__delay_1640__variable_218 <= __delay_data_1640__variable_218;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1644__delay_1643__variable_219 <= __delay_data_1643__variable_219;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1647__delay_1646__variable_220 <= __delay_data_1646__variable_220;
      end 
      if(_mul_10_stream_oready) begin
        _cond_data_231 <= (__delay_data_1637_greaterthan_221)? _sll_data_225 : 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1639__delay_1638_greatereq_234 <= __delay_data_1638_greatereq_234;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1642__delay_1641__delay_1640__variable_218 <= __delay_data_1641__delay_1640__variable_218;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1645__delay_1644__delay_1643__variable_219 <= __delay_data_1644__delay_1643__variable_219;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1648__delay_1647__delay_1646__variable_220 <= __delay_data_1647__delay_1646__variable_220;
      end 
      if(_mul_10_stream_oready) begin
        __muladd_madd_odata_reg_237 <= __muladd_madd_odata_237;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1649__delay_1648__delay_1647____variable_220 <= __delay_data_1648__delay_1647__delay_1646__variable_220;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1650__delay_1649__delay_1648____variable_220 <= __delay_data_1649__delay_1648__delay_1647____variable_220;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1651__delay_1650__delay_1649____variable_220 <= __delay_data_1650__delay_1649__delay_1648____variable_220;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_1652__delay_1651__delay_1650____variable_220 <= __delay_data_1651__delay_1650__delay_1649____variable_220;
      end 
      if(_mul_10_stream_oready) begin
        _sra_data_238 <= __muladd_data_237 >>> __delay_data_1652__delay_1651__delay_1650____variable_220;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_218 <= _cond_data_1585;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_219 <= _cond_data_1423;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_220 <= __delay_data_2698__delay_2697_plus_1653;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_556 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_557 <= _tmp_556;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_558 <= _tmp_557;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_559 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_560 <= _tmp_559;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_561 <= _tmp_560;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_562 <= _tmp_561;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_563 <= _tmp_562;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_564 <= _tmp_563;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_565 <= _tmp_564;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_566 <= _tmp_565;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_567 <= _tmp_566;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_568 <= _tmp_567;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_569 <= _mul_10_source_stop;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_570 <= _tmp_569;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_571 <= _tmp_570;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_572 <= _tmp_571;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_573 <= _tmp_572;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_574 <= _tmp_573;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_575 <= _tmp_574;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_576 <= _tmp_575;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_577 <= _tmp_576;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_578 <= _tmp_577;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_579 <= _mul_10_source_busy;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_580 <= _tmp_579;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_581 <= _tmp_580;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_582 <= _tmp_581;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_583 <= _tmp_582;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_584 <= _tmp_583;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_585 <= _tmp_584;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_586 <= _tmp_585;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_587 <= _tmp_586;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_588 <= _tmp_587;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_589 <= _mul_10_sink_busy;
      end 
      if(!_mul_10_sink_busy && _tmp_589) begin
        _mul_10_busy_reg <= 0;
      end 
      if(_mul_10_source_busy) begin
        _mul_10_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_218 <= _cond_data_2611;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_219 <= _cond_data_2574;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_220 <= __delay_data_3186__delay_3185_plus_2613;
      end 
    end
  end

  localparam _mul_10_fsm_1 = 1;
  localparam _mul_10_fsm_2 = 2;
  localparam _mul_10_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_fsm <= _mul_10_fsm_init;
      _mul_10_source_start <= 0;
      _mul_10_source_busy <= 0;
      _mul_10_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_10_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_10_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_10_stream_oready && _tmp_558) begin
        _mul_10_stream_ivalid <= 1;
      end 
      if(_mul_10_stream_oready && 1'd0) begin
        _mul_10_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        _mul_10_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _mul_10_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_mul_10_fsm)
        _mul_10_fsm_init: begin
          if(_mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
        _mul_10_fsm_1: begin
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_source_start <= 0;
            _mul_10_source_busy <= 1;
          end 
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_2;
          end 
        end
        _mul_10_fsm_2: begin
          if(_mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_3;
          end 
        end
        _mul_10_fsm_3: begin
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_source_busy <= 0;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_fsm <= _mul_10_fsm_init;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_x_source_ram_renable <= 0;
      _mul_11_x_source_fifo_deq <= 0;
      _mul_11_x_idle <= 1;
      _mul_11_y_source_ram_renable <= 0;
      _mul_11_y_source_fifo_deq <= 0;
      _mul_11_y_idle <= 1;
      _mul_11_rshift_source_ram_renable <= 0;
      _mul_11_rshift_source_fifo_deq <= 0;
      _mul_11_rshift_idle <= 1;
      _mul_11_z_sink_wenable <= 0;
      _mul_11_z_sink_fifo_enq <= 0;
      __mul_11_stream_ivalid_1 <= 0;
      __mul_11_stream_ivalid_2 <= 0;
      __mul_11_stream_ivalid_3 <= 0;
      __mul_11_stream_ivalid_4 <= 0;
      __mul_11_stream_ivalid_5 <= 0;
      __mul_11_stream_ivalid_6 <= 0;
      __mul_11_stream_ivalid_7 <= 0;
      __mul_11_stream_ivalid_8 <= 0;
      _greaterthan_data_242 <= 0;
      _minus_data_244 <= 0;
      _greatereq_data_255 <= 0;
      __delay_data_1659__variable_239 <= 0;
      __delay_data_1662__variable_240 <= 0;
      __delay_data_1665__variable_241 <= 0;
      _sll_data_246 <= 0;
      __delay_data_1656_greaterthan_242 <= 0;
      __delay_data_1657_greatereq_255 <= 0;
      __delay_data_1660__delay_1659__variable_239 <= 0;
      __delay_data_1663__delay_1662__variable_240 <= 0;
      __delay_data_1666__delay_1665__variable_241 <= 0;
      _cond_data_252 <= 0;
      __delay_data_1658__delay_1657_greatereq_255 <= 0;
      __delay_data_1661__delay_1660__delay_1659__variable_239 <= 0;
      __delay_data_1664__delay_1663__delay_1662__variable_240 <= 0;
      __delay_data_1667__delay_1666__delay_1665__variable_241 <= 0;
      __muladd_madd_odata_reg_258 <= 0;
      __delay_data_1668__delay_1667__delay_1666____variable_241 <= 0;
      __delay_data_1669__delay_1668__delay_1667____variable_241 <= 0;
      __delay_data_1670__delay_1669__delay_1668____variable_241 <= 0;
      __delay_data_1671__delay_1670__delay_1669____variable_241 <= 0;
      _sra_data_259 <= 0;
      __variable_wdata_239 <= 0;
      __variable_wdata_240 <= 0;
      __variable_wdata_241 <= 0;
      _tmp_590 <= 0;
      _tmp_591 <= 0;
      _tmp_592 <= 0;
      _tmp_593 <= 0;
      _tmp_594 <= 0;
      _tmp_595 <= 0;
      _tmp_596 <= 0;
      _tmp_597 <= 0;
      _tmp_598 <= 0;
      _tmp_599 <= 0;
      _tmp_600 <= 0;
      _tmp_601 <= 0;
      _tmp_602 <= 0;
      _tmp_603 <= 0;
      _tmp_604 <= 0;
      _tmp_605 <= 0;
      _tmp_606 <= 0;
      _tmp_607 <= 0;
      _tmp_608 <= 0;
      _tmp_609 <= 0;
      _tmp_610 <= 0;
      _tmp_611 <= 0;
      _tmp_612 <= 0;
      _tmp_613 <= 0;
      _tmp_614 <= 0;
      _tmp_615 <= 0;
      _tmp_616 <= 0;
      _tmp_617 <= 0;
      _tmp_618 <= 0;
      _tmp_619 <= 0;
      _tmp_620 <= 0;
      _tmp_621 <= 0;
      _tmp_622 <= 0;
      _tmp_623 <= 0;
      _mul_11_busy_reg <= 0;
    end else begin
      if(_mul_11_stream_oready) begin
        _mul_11_x_source_ram_renable <= 0;
        _mul_11_x_source_fifo_deq <= 0;
      end 
      _mul_11_x_idle <= _mul_11_x_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_y_source_ram_renable <= 0;
        _mul_11_y_source_fifo_deq <= 0;
      end 
      _mul_11_y_idle <= _mul_11_y_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_rshift_source_ram_renable <= 0;
        _mul_11_rshift_source_fifo_deq <= 0;
      end 
      _mul_11_rshift_idle <= _mul_11_rshift_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_z_sink_wenable <= 0;
        _mul_11_z_sink_fifo_enq <= 0;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_1 <= _mul_11_stream_ivalid;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_2 <= __mul_11_stream_ivalid_1;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_3 <= __mul_11_stream_ivalid_2;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_4 <= __mul_11_stream_ivalid_3;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_5 <= __mul_11_stream_ivalid_4;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_6 <= __mul_11_stream_ivalid_5;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_7 <= __mul_11_stream_ivalid_6;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_8 <= __mul_11_stream_ivalid_7;
      end 
      if(_mul_11_stream_oready) begin
        _greaterthan_data_242 <= mul_11_rshift_data > 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        _minus_data_244 <= mul_11_rshift_data - 2'sd1;
      end 
      if(_mul_11_stream_oready) begin
        _greatereq_data_255 <= mul_11_x_data >= 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1659__variable_239 <= mul_11_x_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1662__variable_240 <= mul_11_y_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1665__variable_241 <= mul_11_rshift_data;
      end 
      if(_mul_11_stream_oready) begin
        _sll_data_246 <= 2'sd1 << _minus_data_244;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1656_greaterthan_242 <= _greaterthan_data_242;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1657_greatereq_255 <= _greatereq_data_255;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1660__delay_1659__variable_239 <= __delay_data_1659__variable_239;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1663__delay_1662__variable_240 <= __delay_data_1662__variable_240;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1666__delay_1665__variable_241 <= __delay_data_1665__variable_241;
      end 
      if(_mul_11_stream_oready) begin
        _cond_data_252 <= (__delay_data_1656_greaterthan_242)? _sll_data_246 : 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1658__delay_1657_greatereq_255 <= __delay_data_1657_greatereq_255;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1661__delay_1660__delay_1659__variable_239 <= __delay_data_1660__delay_1659__variable_239;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1664__delay_1663__delay_1662__variable_240 <= __delay_data_1663__delay_1662__variable_240;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1667__delay_1666__delay_1665__variable_241 <= __delay_data_1666__delay_1665__variable_241;
      end 
      if(_mul_11_stream_oready) begin
        __muladd_madd_odata_reg_258 <= __muladd_madd_odata_258;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1668__delay_1667__delay_1666____variable_241 <= __delay_data_1667__delay_1666__delay_1665__variable_241;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1669__delay_1668__delay_1667____variable_241 <= __delay_data_1668__delay_1667__delay_1666____variable_241;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1670__delay_1669__delay_1668____variable_241 <= __delay_data_1669__delay_1668__delay_1667____variable_241;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_1671__delay_1670__delay_1669____variable_241 <= __delay_data_1670__delay_1669__delay_1668____variable_241;
      end 
      if(_mul_11_stream_oready) begin
        _sra_data_259 <= __muladd_data_258 >>> __delay_data_1671__delay_1670__delay_1669____variable_241;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_239 <= _cond_data_1587;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_240 <= _cond_data_1425;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_241 <= __delay_data_2715__delay_2714_plus_1672;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_590 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_591 <= _tmp_590;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_592 <= _tmp_591;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_593 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_594 <= _tmp_593;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_595 <= _tmp_594;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_596 <= _tmp_595;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_597 <= _tmp_596;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_598 <= _tmp_597;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_599 <= _tmp_598;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_600 <= _tmp_599;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_601 <= _tmp_600;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_602 <= _tmp_601;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_603 <= _mul_11_source_stop;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_604 <= _tmp_603;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_605 <= _tmp_604;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_606 <= _tmp_605;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_607 <= _tmp_606;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_608 <= _tmp_607;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_609 <= _tmp_608;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_610 <= _tmp_609;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_611 <= _tmp_610;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_612 <= _tmp_611;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_613 <= _mul_11_source_busy;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_614 <= _tmp_613;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_615 <= _tmp_614;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_616 <= _tmp_615;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_617 <= _tmp_616;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_618 <= _tmp_617;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_619 <= _tmp_618;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_620 <= _tmp_619;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_621 <= _tmp_620;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_622 <= _tmp_621;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_623 <= _mul_11_sink_busy;
      end 
      if(!_mul_11_sink_busy && _tmp_623) begin
        _mul_11_busy_reg <= 0;
      end 
      if(_mul_11_source_busy) begin
        _mul_11_busy_reg <= 1;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_239 <= _cond_data_2616;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_240 <= _cond_data_2576;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        __variable_wdata_241 <= __delay_data_3191__delay_3190_plus_2618;
      end 
    end
  end

  localparam _mul_11_fsm_1 = 1;
  localparam _mul_11_fsm_2 = 2;
  localparam _mul_11_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_fsm <= _mul_11_fsm_init;
      _mul_11_source_start <= 0;
      _mul_11_source_busy <= 0;
      _mul_11_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_11_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_11_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_11_stream_oready && _tmp_592) begin
        _mul_11_stream_ivalid <= 1;
      end 
      if(_mul_11_stream_oready && 1'd0) begin
        _mul_11_stream_ivalid <= 0;
      end 
      if(__stream_matmul_16_stream_ivalid_3 && _stream_matmul_16_stream_oready) begin
        _mul_11_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_busy) begin
        _mul_11_source_busy <= _stream_matmul_16_source_busy;
      end 
      case(_mul_11_fsm)
        _mul_11_fsm_init: begin
          if(_mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
        _mul_11_fsm_1: begin
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_source_start <= 0;
            _mul_11_source_busy <= 1;
          end 
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_2;
          end 
        end
        _mul_11_fsm_2: begin
          if(_mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_3;
          end 
        end
        _mul_11_fsm_3: begin
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_source_busy <= 0;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_fsm <= _mul_11_fsm_init;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_x_source_ram_renable <= 0;
      _mul_12_x_source_fifo_deq <= 0;
      _mul_12_x_idle <= 1;
      _mul_12_y_source_ram_renable <= 0;
      _mul_12_y_source_fifo_deq <= 0;
      _mul_12_y_idle <= 1;
      _mul_12_rshift_source_ram_renable <= 0;
      _mul_12_rshift_source_fifo_deq <= 0;
      _mul_12_rshift_idle <= 1;
      _mul_12_z_sink_wenable <= 0;
      _mul_12_z_sink_fifo_enq <= 0;
      __mul_12_stream_ivalid_1 <= 0;
      __mul_12_stream_ivalid_2 <= 0;
      __mul_12_stream_ivalid_3 <= 0;
      __mul_12_stream_ivalid_4 <= 0;
      __mul_12_stream_ivalid_5 <= 0;
      __mul_12_stream_ivalid_6 <= 0;
      __mul_12_stream_ivalid_7 <= 0;
      __mul_12_stream_ivalid_8 <= 0;
      _greaterthan_data_263 <= 0;
      _minus_data_265 <= 0;
      _greatereq_data_276 <= 0;
      __delay_data_1678__variable_260 <= 0;
      __delay_data_1681__variable_261 <= 0;
      __delay_data_1684__variable_262 <= 0;
      _sll_data_267 <= 0;
      __delay_data_1675_greaterthan_263 <= 0;
      __delay_data_1676_greatereq_276 <= 0;
      __delay_data_1679__delay_1678__variable_260 <= 0;
      __delay_data_1682__delay_1681__variable_261 <= 0;
      __delay_data_1685__delay_1684__variable_262 <= 0;
      _cond_data_273 <= 0;
      __delay_data_1677__delay_1676_greatereq_276 <= 0;
      __delay_data_1680__delay_1679__delay_1678__variable_260 <= 0;
      __delay_data_1683__delay_1682__delay_1681__variable_261 <= 0;
      __delay_data_1686__delay_1685__delay_1684__variable_262 <= 0;
      __muladd_madd_odata_reg_279 <= 0;
      __delay_data_1687__delay_1686__delay_1685____variable_262 <= 0;
      __delay_data_1688__delay_1687__delay_1686____variable_262 <= 0;
      __delay_data_1689__delay_1688__delay_1687____variable_262 <= 0;
      __delay_data_1690__delay_1689__delay_1688____variable_262 <= 0;
      _sra_data_280 <= 0;
      __variable_wdata_260 <= 0;
      __variable_wdata_261 <= 0;
      __variable_wdata_262 <= 0;
      _tmp_624 <= 0;
      _tmp_625 <= 0;
      _tmp_626 <= 0;
      _tmp_627 <= 0;
      _tmp_628 <= 0;
      _tmp_629 <= 0;
      _tmp_630 <= 0;
      _tmp_631 <= 0;
      _tmp_632 <= 0;
      _tmp_633 <= 0;
      _tmp_634 <= 0;
      _tmp_635 <= 0;
      _tmp_636 <= 0;
      _tmp_637 <= 0;
      _tmp_638 <= 0;
      _tmp_639 <= 0;
      _tmp_640 <= 0;
      _tmp_641 <= 0;
      _tmp_642 <= 0;
      _tmp_643 <= 0;
      _tmp_644 <= 0;
      _tmp_645 <= 0;
      _tmp_646 <= 0;
      _tmp_647 <= 0;
      _tmp_648 <= 0;
      _tmp_649 <= 0;
      _tmp_650 <= 0;
      _tmp_651 <= 0;
      _tmp_652 <= 0;
      _tmp_653 <= 0;
      _tmp_654 <= 0;
      _tmp_655 <= 0;
      _tmp_656 <= 0;
      _tmp_657 <= 0;
      _mul_12_busy_reg <= 0;
    end else begin
      if(_mul_12_stream_oready) begin
        _mul_12_x_source_ram_renable <= 0;
        _mul_12_x_source_fifo_deq <= 0;
      end 
      _mul_12_x_idle <= _mul_12_x_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_y_source_ram_renable <= 0;
        _mul_12_y_source_fifo_deq <= 0;
      end 
      _mul_12_y_idle <= _mul_12_y_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_rshift_source_ram_renable <= 0;
        _mul_12_rshift_source_fifo_deq <= 0;
      end 
      _mul_12_rshift_idle <= _mul_12_rshift_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_z_sink_wenable <= 0;
        _mul_12_z_sink_fifo_enq <= 0;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_1 <= _mul_12_stream_ivalid;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_2 <= __mul_12_stream_ivalid_1;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_3 <= __mul_12_stream_ivalid_2;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_4 <= __mul_12_stream_ivalid_3;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_5 <= __mul_12_stream_ivalid_4;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_6 <= __mul_12_stream_ivalid_5;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_7 <= __mul_12_stream_ivalid_6;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_8 <= __mul_12_stream_ivalid_7;
      end 
      if(_mul_12_stream_oready) begin
        _greaterthan_data_263 <= mul_12_rshift_data > 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        _minus_data_265 <= mul_12_rshift_data - 2'sd1;
      end 
      if(_mul_12_stream_oready) begin
        _greatereq_data_276 <= mul_12_x_data >= 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1678__variable_260 <= mul_12_x_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1681__variable_261 <= mul_12_y_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1684__variable_262 <= mul_12_rshift_data;
      end 
      if(_mul_12_stream_oready) begin
        _sll_data_267 <= 2'sd1 << _minus_data_265;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1675_greaterthan_263 <= _greaterthan_data_263;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1676_greatereq_276 <= _greatereq_data_276;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1679__delay_1678__variable_260 <= __delay_data_1678__variable_260;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1682__delay_1681__variable_261 <= __delay_data_1681__variable_261;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1685__delay_1684__variable_262 <= __delay_data_1684__variable_262;
      end 
      if(_mul_12_stream_oready) begin
        _cond_data_273 <= (__delay_data_1675_greaterthan_263)? _sll_data_267 : 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1677__delay_1676_greatereq_276 <= __delay_data_1676_greatereq_276;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1680__delay_1679__delay_1678__variable_260 <= __delay_data_1679__delay_1678__variable_260;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1683__delay_1682__delay_1681__variable_261 <= __delay_data_1682__delay_1681__variable_261;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1686__delay_1685__delay_1684__variable_262 <= __delay_data_1685__delay_1684__variable_262;
      end 
      if(_mul_12_stream_oready) begin
        __muladd_madd_odata_reg_279 <= __muladd_madd_odata_279;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1687__delay_1686__delay_1685____variable_262 <= __delay_data_1686__delay_1685__delay_1684__variable_262;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1688__delay_1687__delay_1686____variable_262 <= __delay_data_1687__delay_1686__delay_1685____variable_262;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1689__delay_1688__delay_1687____variable_262 <= __delay_data_1688__delay_1687__delay_1686____variable_262;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_1690__delay_1689__delay_1688____variable_262 <= __delay_data_1689__delay_1688__delay_1687____variable_262;
      end 
      if(_mul_12_stream_oready) begin
        _sra_data_280 <= __muladd_data_279 >>> __delay_data_1690__delay_1689__delay_1688____variable_262;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_260 <= _cond_data_1589;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_261 <= _cond_data_1427;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_262 <= __delay_data_2732__delay_2731_plus_1691;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_624 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_625 <= _tmp_624;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_626 <= _tmp_625;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_627 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_628 <= _tmp_627;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_629 <= _tmp_628;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_630 <= _tmp_629;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_631 <= _tmp_630;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_632 <= _tmp_631;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_633 <= _tmp_632;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_634 <= _tmp_633;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_635 <= _tmp_634;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_636 <= _tmp_635;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_637 <= _mul_12_source_stop;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_638 <= _tmp_637;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_639 <= _tmp_638;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_640 <= _tmp_639;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_641 <= _tmp_640;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_642 <= _tmp_641;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_643 <= _tmp_642;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_644 <= _tmp_643;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_645 <= _tmp_644;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_646 <= _tmp_645;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_647 <= _mul_12_source_busy;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_648 <= _tmp_647;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_649 <= _tmp_648;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_650 <= _tmp_649;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_651 <= _tmp_650;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_652 <= _tmp_651;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_653 <= _tmp_652;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_654 <= _tmp_653;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_655 <= _tmp_654;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_656 <= _tmp_655;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_657 <= _mul_12_sink_busy;
      end 
      if(!_mul_12_sink_busy && _tmp_657) begin
        _mul_12_busy_reg <= 0;
      end 
      if(_mul_12_source_busy) begin
        _mul_12_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_12_fsm_1 = 1;
  localparam _mul_12_fsm_2 = 2;
  localparam _mul_12_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_fsm <= _mul_12_fsm_init;
      _mul_12_source_start <= 0;
      _mul_12_source_busy <= 0;
      _mul_12_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_12_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_12_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_12_stream_oready && _tmp_626) begin
        _mul_12_stream_ivalid <= 1;
      end 
      if(_mul_12_stream_oready && 1'd0) begin
        _mul_12_stream_ivalid <= 0;
      end 
      case(_mul_12_fsm)
        _mul_12_fsm_init: begin
          if(_mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
        _mul_12_fsm_1: begin
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_source_start <= 0;
            _mul_12_source_busy <= 1;
          end 
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_2;
          end 
        end
        _mul_12_fsm_2: begin
          if(_mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_3;
          end 
        end
        _mul_12_fsm_3: begin
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_source_busy <= 0;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_fsm <= _mul_12_fsm_init;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_13_x_source_ram_renable <= 0;
      _mul_13_x_source_fifo_deq <= 0;
      _mul_13_x_idle <= 1;
      _mul_13_y_source_ram_renable <= 0;
      _mul_13_y_source_fifo_deq <= 0;
      _mul_13_y_idle <= 1;
      _mul_13_rshift_source_ram_renable <= 0;
      _mul_13_rshift_source_fifo_deq <= 0;
      _mul_13_rshift_idle <= 1;
      _mul_13_z_sink_wenable <= 0;
      _mul_13_z_sink_fifo_enq <= 0;
      __mul_13_stream_ivalid_1 <= 0;
      __mul_13_stream_ivalid_2 <= 0;
      __mul_13_stream_ivalid_3 <= 0;
      __mul_13_stream_ivalid_4 <= 0;
      __mul_13_stream_ivalid_5 <= 0;
      __mul_13_stream_ivalid_6 <= 0;
      __mul_13_stream_ivalid_7 <= 0;
      __mul_13_stream_ivalid_8 <= 0;
      _greaterthan_data_284 <= 0;
      _minus_data_286 <= 0;
      _greatereq_data_297 <= 0;
      __delay_data_1697__variable_281 <= 0;
      __delay_data_1700__variable_282 <= 0;
      __delay_data_1703__variable_283 <= 0;
      _sll_data_288 <= 0;
      __delay_data_1694_greaterthan_284 <= 0;
      __delay_data_1695_greatereq_297 <= 0;
      __delay_data_1698__delay_1697__variable_281 <= 0;
      __delay_data_1701__delay_1700__variable_282 <= 0;
      __delay_data_1704__delay_1703__variable_283 <= 0;
      _cond_data_294 <= 0;
      __delay_data_1696__delay_1695_greatereq_297 <= 0;
      __delay_data_1699__delay_1698__delay_1697__variable_281 <= 0;
      __delay_data_1702__delay_1701__delay_1700__variable_282 <= 0;
      __delay_data_1705__delay_1704__delay_1703__variable_283 <= 0;
      __muladd_madd_odata_reg_300 <= 0;
      __delay_data_1706__delay_1705__delay_1704____variable_283 <= 0;
      __delay_data_1707__delay_1706__delay_1705____variable_283 <= 0;
      __delay_data_1708__delay_1707__delay_1706____variable_283 <= 0;
      __delay_data_1709__delay_1708__delay_1707____variable_283 <= 0;
      _sra_data_301 <= 0;
      __variable_wdata_281 <= 0;
      __variable_wdata_282 <= 0;
      __variable_wdata_283 <= 0;
      _tmp_658 <= 0;
      _tmp_659 <= 0;
      _tmp_660 <= 0;
      _tmp_661 <= 0;
      _tmp_662 <= 0;
      _tmp_663 <= 0;
      _tmp_664 <= 0;
      _tmp_665 <= 0;
      _tmp_666 <= 0;
      _tmp_667 <= 0;
      _tmp_668 <= 0;
      _tmp_669 <= 0;
      _tmp_670 <= 0;
      _tmp_671 <= 0;
      _tmp_672 <= 0;
      _tmp_673 <= 0;
      _tmp_674 <= 0;
      _tmp_675 <= 0;
      _tmp_676 <= 0;
      _tmp_677 <= 0;
      _tmp_678 <= 0;
      _tmp_679 <= 0;
      _tmp_680 <= 0;
      _tmp_681 <= 0;
      _tmp_682 <= 0;
      _tmp_683 <= 0;
      _tmp_684 <= 0;
      _tmp_685 <= 0;
      _tmp_686 <= 0;
      _tmp_687 <= 0;
      _tmp_688 <= 0;
      _tmp_689 <= 0;
      _tmp_690 <= 0;
      _tmp_691 <= 0;
      _mul_13_busy_reg <= 0;
    end else begin
      if(_mul_13_stream_oready) begin
        _mul_13_x_source_ram_renable <= 0;
        _mul_13_x_source_fifo_deq <= 0;
      end 
      _mul_13_x_idle <= _mul_13_x_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_y_source_ram_renable <= 0;
        _mul_13_y_source_fifo_deq <= 0;
      end 
      _mul_13_y_idle <= _mul_13_y_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_rshift_source_ram_renable <= 0;
        _mul_13_rshift_source_fifo_deq <= 0;
      end 
      _mul_13_rshift_idle <= _mul_13_rshift_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_z_sink_wenable <= 0;
        _mul_13_z_sink_fifo_enq <= 0;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_1 <= _mul_13_stream_ivalid;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_2 <= __mul_13_stream_ivalid_1;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_3 <= __mul_13_stream_ivalid_2;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_4 <= __mul_13_stream_ivalid_3;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_5 <= __mul_13_stream_ivalid_4;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_6 <= __mul_13_stream_ivalid_5;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_7 <= __mul_13_stream_ivalid_6;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_8 <= __mul_13_stream_ivalid_7;
      end 
      if(_mul_13_stream_oready) begin
        _greaterthan_data_284 <= mul_13_rshift_data > 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        _minus_data_286 <= mul_13_rshift_data - 2'sd1;
      end 
      if(_mul_13_stream_oready) begin
        _greatereq_data_297 <= mul_13_x_data >= 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1697__variable_281 <= mul_13_x_data;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1700__variable_282 <= mul_13_y_data;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1703__variable_283 <= mul_13_rshift_data;
      end 
      if(_mul_13_stream_oready) begin
        _sll_data_288 <= 2'sd1 << _minus_data_286;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1694_greaterthan_284 <= _greaterthan_data_284;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1695_greatereq_297 <= _greatereq_data_297;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1698__delay_1697__variable_281 <= __delay_data_1697__variable_281;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1701__delay_1700__variable_282 <= __delay_data_1700__variable_282;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1704__delay_1703__variable_283 <= __delay_data_1703__variable_283;
      end 
      if(_mul_13_stream_oready) begin
        _cond_data_294 <= (__delay_data_1694_greaterthan_284)? _sll_data_288 : 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1696__delay_1695_greatereq_297 <= __delay_data_1695_greatereq_297;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1699__delay_1698__delay_1697__variable_281 <= __delay_data_1698__delay_1697__variable_281;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1702__delay_1701__delay_1700__variable_282 <= __delay_data_1701__delay_1700__variable_282;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1705__delay_1704__delay_1703__variable_283 <= __delay_data_1704__delay_1703__variable_283;
      end 
      if(_mul_13_stream_oready) begin
        __muladd_madd_odata_reg_300 <= __muladd_madd_odata_300;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1706__delay_1705__delay_1704____variable_283 <= __delay_data_1705__delay_1704__delay_1703__variable_283;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1707__delay_1706__delay_1705____variable_283 <= __delay_data_1706__delay_1705__delay_1704____variable_283;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1708__delay_1707__delay_1706____variable_283 <= __delay_data_1707__delay_1706__delay_1705____variable_283;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_1709__delay_1708__delay_1707____variable_283 <= __delay_data_1708__delay_1707__delay_1706____variable_283;
      end 
      if(_mul_13_stream_oready) begin
        _sra_data_301 <= __muladd_data_300 >>> __delay_data_1709__delay_1708__delay_1707____variable_283;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_281 <= _cond_data_1591;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_282 <= _cond_data_1429;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_283 <= __delay_data_2749__delay_2748_plus_1710;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_658 <= _mul_13_source_start;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_659 <= _tmp_658;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_660 <= _tmp_659;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_661 <= _mul_13_source_start;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_662 <= _tmp_661;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_663 <= _tmp_662;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_664 <= _tmp_663;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_665 <= _tmp_664;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_666 <= _tmp_665;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_667 <= _tmp_666;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_668 <= _tmp_667;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_669 <= _tmp_668;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_670 <= _tmp_669;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_671 <= _mul_13_source_stop;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_672 <= _tmp_671;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_673 <= _tmp_672;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_674 <= _tmp_673;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_675 <= _tmp_674;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_676 <= _tmp_675;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_677 <= _tmp_676;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_678 <= _tmp_677;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_679 <= _tmp_678;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_680 <= _tmp_679;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_681 <= _mul_13_source_busy;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_682 <= _tmp_681;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_683 <= _tmp_682;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_684 <= _tmp_683;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_685 <= _tmp_684;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_686 <= _tmp_685;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_687 <= _tmp_686;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_688 <= _tmp_687;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_689 <= _tmp_688;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_690 <= _tmp_689;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_691 <= _mul_13_sink_busy;
      end 
      if(!_mul_13_sink_busy && _tmp_691) begin
        _mul_13_busy_reg <= 0;
      end 
      if(_mul_13_source_busy) begin
        _mul_13_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_13_fsm_1 = 1;
  localparam _mul_13_fsm_2 = 2;
  localparam _mul_13_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_13_fsm <= _mul_13_fsm_init;
      _mul_13_source_start <= 0;
      _mul_13_source_busy <= 0;
      _mul_13_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_13_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_13_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_13_stream_oready && _tmp_660) begin
        _mul_13_stream_ivalid <= 1;
      end 
      if(_mul_13_stream_oready && 1'd0) begin
        _mul_13_stream_ivalid <= 0;
      end 
      case(_mul_13_fsm)
        _mul_13_fsm_init: begin
          if(_mul_13_run_flag) begin
            _mul_13_source_start <= 1;
          end 
          if(_mul_13_run_flag) begin
            _mul_13_fsm <= _mul_13_fsm_1;
          end 
        end
        _mul_13_fsm_1: begin
          if(_mul_13_source_start && _mul_13_stream_oready) begin
            _mul_13_source_start <= 0;
            _mul_13_source_busy <= 1;
          end 
          if(_mul_13_source_start && _mul_13_stream_oready) begin
            _mul_13_fsm <= _mul_13_fsm_2;
          end 
        end
        _mul_13_fsm_2: begin
          if(_mul_13_stream_oready) begin
            _mul_13_fsm <= _mul_13_fsm_3;
          end 
        end
        _mul_13_fsm_3: begin
          if(_mul_13_stream_oready && 1'd0) begin
            _mul_13_source_busy <= 0;
          end 
          if(_mul_13_stream_oready && 1'd0 && _mul_13_run_flag) begin
            _mul_13_source_start <= 1;
          end 
          if(_mul_13_stream_oready && 1'd0) begin
            _mul_13_fsm <= _mul_13_fsm_init;
          end 
          if(_mul_13_stream_oready && 1'd0 && _mul_13_run_flag) begin
            _mul_13_fsm <= _mul_13_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_14_x_source_ram_renable <= 0;
      _mul_14_x_source_fifo_deq <= 0;
      _mul_14_x_idle <= 1;
      _mul_14_y_source_ram_renable <= 0;
      _mul_14_y_source_fifo_deq <= 0;
      _mul_14_y_idle <= 1;
      _mul_14_rshift_source_ram_renable <= 0;
      _mul_14_rshift_source_fifo_deq <= 0;
      _mul_14_rshift_idle <= 1;
      _mul_14_z_sink_wenable <= 0;
      _mul_14_z_sink_fifo_enq <= 0;
      __mul_14_stream_ivalid_1 <= 0;
      __mul_14_stream_ivalid_2 <= 0;
      __mul_14_stream_ivalid_3 <= 0;
      __mul_14_stream_ivalid_4 <= 0;
      __mul_14_stream_ivalid_5 <= 0;
      __mul_14_stream_ivalid_6 <= 0;
      __mul_14_stream_ivalid_7 <= 0;
      __mul_14_stream_ivalid_8 <= 0;
      _greaterthan_data_305 <= 0;
      _minus_data_307 <= 0;
      _greatereq_data_318 <= 0;
      __delay_data_1716__variable_302 <= 0;
      __delay_data_1719__variable_303 <= 0;
      __delay_data_1722__variable_304 <= 0;
      _sll_data_309 <= 0;
      __delay_data_1713_greaterthan_305 <= 0;
      __delay_data_1714_greatereq_318 <= 0;
      __delay_data_1717__delay_1716__variable_302 <= 0;
      __delay_data_1720__delay_1719__variable_303 <= 0;
      __delay_data_1723__delay_1722__variable_304 <= 0;
      _cond_data_315 <= 0;
      __delay_data_1715__delay_1714_greatereq_318 <= 0;
      __delay_data_1718__delay_1717__delay_1716__variable_302 <= 0;
      __delay_data_1721__delay_1720__delay_1719__variable_303 <= 0;
      __delay_data_1724__delay_1723__delay_1722__variable_304 <= 0;
      __muladd_madd_odata_reg_321 <= 0;
      __delay_data_1725__delay_1724__delay_1723____variable_304 <= 0;
      __delay_data_1726__delay_1725__delay_1724____variable_304 <= 0;
      __delay_data_1727__delay_1726__delay_1725____variable_304 <= 0;
      __delay_data_1728__delay_1727__delay_1726____variable_304 <= 0;
      _sra_data_322 <= 0;
      __variable_wdata_302 <= 0;
      __variable_wdata_303 <= 0;
      __variable_wdata_304 <= 0;
      _tmp_692 <= 0;
      _tmp_693 <= 0;
      _tmp_694 <= 0;
      _tmp_695 <= 0;
      _tmp_696 <= 0;
      _tmp_697 <= 0;
      _tmp_698 <= 0;
      _tmp_699 <= 0;
      _tmp_700 <= 0;
      _tmp_701 <= 0;
      _tmp_702 <= 0;
      _tmp_703 <= 0;
      _tmp_704 <= 0;
      _tmp_705 <= 0;
      _tmp_706 <= 0;
      _tmp_707 <= 0;
      _tmp_708 <= 0;
      _tmp_709 <= 0;
      _tmp_710 <= 0;
      _tmp_711 <= 0;
      _tmp_712 <= 0;
      _tmp_713 <= 0;
      _tmp_714 <= 0;
      _tmp_715 <= 0;
      _tmp_716 <= 0;
      _tmp_717 <= 0;
      _tmp_718 <= 0;
      _tmp_719 <= 0;
      _tmp_720 <= 0;
      _tmp_721 <= 0;
      _tmp_722 <= 0;
      _tmp_723 <= 0;
      _tmp_724 <= 0;
      _tmp_725 <= 0;
      _mul_14_busy_reg <= 0;
    end else begin
      if(_mul_14_stream_oready) begin
        _mul_14_x_source_ram_renable <= 0;
        _mul_14_x_source_fifo_deq <= 0;
      end 
      _mul_14_x_idle <= _mul_14_x_idle;
      if(_mul_14_stream_oready) begin
        _mul_14_y_source_ram_renable <= 0;
        _mul_14_y_source_fifo_deq <= 0;
      end 
      _mul_14_y_idle <= _mul_14_y_idle;
      if(_mul_14_stream_oready) begin
        _mul_14_rshift_source_ram_renable <= 0;
        _mul_14_rshift_source_fifo_deq <= 0;
      end 
      _mul_14_rshift_idle <= _mul_14_rshift_idle;
      if(_mul_14_stream_oready) begin
        _mul_14_z_sink_wenable <= 0;
        _mul_14_z_sink_fifo_enq <= 0;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_1 <= _mul_14_stream_ivalid;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_2 <= __mul_14_stream_ivalid_1;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_3 <= __mul_14_stream_ivalid_2;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_4 <= __mul_14_stream_ivalid_3;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_5 <= __mul_14_stream_ivalid_4;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_6 <= __mul_14_stream_ivalid_5;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_7 <= __mul_14_stream_ivalid_6;
      end 
      if(_mul_14_stream_oready) begin
        __mul_14_stream_ivalid_8 <= __mul_14_stream_ivalid_7;
      end 
      if(_mul_14_stream_oready) begin
        _greaterthan_data_305 <= mul_14_rshift_data > 1'sd0;
      end 
      if(_mul_14_stream_oready) begin
        _minus_data_307 <= mul_14_rshift_data - 2'sd1;
      end 
      if(_mul_14_stream_oready) begin
        _greatereq_data_318 <= mul_14_x_data >= 1'sd0;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1716__variable_302 <= mul_14_x_data;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1719__variable_303 <= mul_14_y_data;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1722__variable_304 <= mul_14_rshift_data;
      end 
      if(_mul_14_stream_oready) begin
        _sll_data_309 <= 2'sd1 << _minus_data_307;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1713_greaterthan_305 <= _greaterthan_data_305;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1714_greatereq_318 <= _greatereq_data_318;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1717__delay_1716__variable_302 <= __delay_data_1716__variable_302;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1720__delay_1719__variable_303 <= __delay_data_1719__variable_303;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1723__delay_1722__variable_304 <= __delay_data_1722__variable_304;
      end 
      if(_mul_14_stream_oready) begin
        _cond_data_315 <= (__delay_data_1713_greaterthan_305)? _sll_data_309 : 1'sd0;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1715__delay_1714_greatereq_318 <= __delay_data_1714_greatereq_318;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1718__delay_1717__delay_1716__variable_302 <= __delay_data_1717__delay_1716__variable_302;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1721__delay_1720__delay_1719__variable_303 <= __delay_data_1720__delay_1719__variable_303;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1724__delay_1723__delay_1722__variable_304 <= __delay_data_1723__delay_1722__variable_304;
      end 
      if(_mul_14_stream_oready) begin
        __muladd_madd_odata_reg_321 <= __muladd_madd_odata_321;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1725__delay_1724__delay_1723____variable_304 <= __delay_data_1724__delay_1723__delay_1722__variable_304;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1726__delay_1725__delay_1724____variable_304 <= __delay_data_1725__delay_1724__delay_1723____variable_304;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1727__delay_1726__delay_1725____variable_304 <= __delay_data_1726__delay_1725__delay_1724____variable_304;
      end 
      if(_mul_14_stream_oready) begin
        __delay_data_1728__delay_1727__delay_1726____variable_304 <= __delay_data_1727__delay_1726__delay_1725____variable_304;
      end 
      if(_mul_14_stream_oready) begin
        _sra_data_322 <= __muladd_data_321 >>> __delay_data_1728__delay_1727__delay_1726____variable_304;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_302 <= _cond_data_1593;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_303 <= _cond_data_1431;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_304 <= __delay_data_2766__delay_2765_plus_1729;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_692 <= _mul_14_source_start;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_693 <= _tmp_692;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_694 <= _tmp_693;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_695 <= _mul_14_source_start;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_696 <= _tmp_695;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_697 <= _tmp_696;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_698 <= _tmp_697;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_699 <= _tmp_698;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_700 <= _tmp_699;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_701 <= _tmp_700;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_702 <= _tmp_701;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_703 <= _tmp_702;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_704 <= _tmp_703;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_705 <= _mul_14_source_stop;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_706 <= _tmp_705;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_707 <= _tmp_706;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_708 <= _tmp_707;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_709 <= _tmp_708;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_710 <= _tmp_709;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_711 <= _tmp_710;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_712 <= _tmp_711;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_713 <= _tmp_712;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_714 <= _tmp_713;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_715 <= _mul_14_source_busy;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_716 <= _tmp_715;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_717 <= _tmp_716;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_718 <= _tmp_717;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_719 <= _tmp_718;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_720 <= _tmp_719;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_721 <= _tmp_720;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_722 <= _tmp_721;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_723 <= _tmp_722;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_724 <= _tmp_723;
      end 
      if(_mul_14_stream_oready) begin
        _tmp_725 <= _mul_14_sink_busy;
      end 
      if(!_mul_14_sink_busy && _tmp_725) begin
        _mul_14_busy_reg <= 0;
      end 
      if(_mul_14_source_busy) begin
        _mul_14_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_14_fsm_1 = 1;
  localparam _mul_14_fsm_2 = 2;
  localparam _mul_14_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_14_fsm <= _mul_14_fsm_init;
      _mul_14_source_start <= 0;
      _mul_14_source_busy <= 0;
      _mul_14_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_14_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_14_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_14_stream_oready && _tmp_694) begin
        _mul_14_stream_ivalid <= 1;
      end 
      if(_mul_14_stream_oready && 1'd0) begin
        _mul_14_stream_ivalid <= 0;
      end 
      case(_mul_14_fsm)
        _mul_14_fsm_init: begin
          if(_mul_14_run_flag) begin
            _mul_14_source_start <= 1;
          end 
          if(_mul_14_run_flag) begin
            _mul_14_fsm <= _mul_14_fsm_1;
          end 
        end
        _mul_14_fsm_1: begin
          if(_mul_14_source_start && _mul_14_stream_oready) begin
            _mul_14_source_start <= 0;
            _mul_14_source_busy <= 1;
          end 
          if(_mul_14_source_start && _mul_14_stream_oready) begin
            _mul_14_fsm <= _mul_14_fsm_2;
          end 
        end
        _mul_14_fsm_2: begin
          if(_mul_14_stream_oready) begin
            _mul_14_fsm <= _mul_14_fsm_3;
          end 
        end
        _mul_14_fsm_3: begin
          if(_mul_14_stream_oready && 1'd0) begin
            _mul_14_source_busy <= 0;
          end 
          if(_mul_14_stream_oready && 1'd0 && _mul_14_run_flag) begin
            _mul_14_source_start <= 1;
          end 
          if(_mul_14_stream_oready && 1'd0) begin
            _mul_14_fsm <= _mul_14_fsm_init;
          end 
          if(_mul_14_stream_oready && 1'd0 && _mul_14_run_flag) begin
            _mul_14_fsm <= _mul_14_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_15_x_source_ram_renable <= 0;
      _mul_15_x_source_fifo_deq <= 0;
      _mul_15_x_idle <= 1;
      _mul_15_y_source_ram_renable <= 0;
      _mul_15_y_source_fifo_deq <= 0;
      _mul_15_y_idle <= 1;
      _mul_15_rshift_source_ram_renable <= 0;
      _mul_15_rshift_source_fifo_deq <= 0;
      _mul_15_rshift_idle <= 1;
      _mul_15_z_sink_wenable <= 0;
      _mul_15_z_sink_fifo_enq <= 0;
      __mul_15_stream_ivalid_1 <= 0;
      __mul_15_stream_ivalid_2 <= 0;
      __mul_15_stream_ivalid_3 <= 0;
      __mul_15_stream_ivalid_4 <= 0;
      __mul_15_stream_ivalid_5 <= 0;
      __mul_15_stream_ivalid_6 <= 0;
      __mul_15_stream_ivalid_7 <= 0;
      __mul_15_stream_ivalid_8 <= 0;
      _greaterthan_data_326 <= 0;
      _minus_data_328 <= 0;
      _greatereq_data_339 <= 0;
      __delay_data_1735__variable_323 <= 0;
      __delay_data_1738__variable_324 <= 0;
      __delay_data_1741__variable_325 <= 0;
      _sll_data_330 <= 0;
      __delay_data_1732_greaterthan_326 <= 0;
      __delay_data_1733_greatereq_339 <= 0;
      __delay_data_1736__delay_1735__variable_323 <= 0;
      __delay_data_1739__delay_1738__variable_324 <= 0;
      __delay_data_1742__delay_1741__variable_325 <= 0;
      _cond_data_336 <= 0;
      __delay_data_1734__delay_1733_greatereq_339 <= 0;
      __delay_data_1737__delay_1736__delay_1735__variable_323 <= 0;
      __delay_data_1740__delay_1739__delay_1738__variable_324 <= 0;
      __delay_data_1743__delay_1742__delay_1741__variable_325 <= 0;
      __muladd_madd_odata_reg_342 <= 0;
      __delay_data_1744__delay_1743__delay_1742____variable_325 <= 0;
      __delay_data_1745__delay_1744__delay_1743____variable_325 <= 0;
      __delay_data_1746__delay_1745__delay_1744____variable_325 <= 0;
      __delay_data_1747__delay_1746__delay_1745____variable_325 <= 0;
      _sra_data_343 <= 0;
      __variable_wdata_323 <= 0;
      __variable_wdata_324 <= 0;
      __variable_wdata_325 <= 0;
      _tmp_726 <= 0;
      _tmp_727 <= 0;
      _tmp_728 <= 0;
      _tmp_729 <= 0;
      _tmp_730 <= 0;
      _tmp_731 <= 0;
      _tmp_732 <= 0;
      _tmp_733 <= 0;
      _tmp_734 <= 0;
      _tmp_735 <= 0;
      _tmp_736 <= 0;
      _tmp_737 <= 0;
      _tmp_738 <= 0;
      _tmp_739 <= 0;
      _tmp_740 <= 0;
      _tmp_741 <= 0;
      _tmp_742 <= 0;
      _tmp_743 <= 0;
      _tmp_744 <= 0;
      _tmp_745 <= 0;
      _tmp_746 <= 0;
      _tmp_747 <= 0;
      _tmp_748 <= 0;
      _tmp_749 <= 0;
      _tmp_750 <= 0;
      _tmp_751 <= 0;
      _tmp_752 <= 0;
      _tmp_753 <= 0;
      _tmp_754 <= 0;
      _tmp_755 <= 0;
      _tmp_756 <= 0;
      _tmp_757 <= 0;
      _tmp_758 <= 0;
      _tmp_759 <= 0;
      _mul_15_busy_reg <= 0;
    end else begin
      if(_mul_15_stream_oready) begin
        _mul_15_x_source_ram_renable <= 0;
        _mul_15_x_source_fifo_deq <= 0;
      end 
      _mul_15_x_idle <= _mul_15_x_idle;
      if(_mul_15_stream_oready) begin
        _mul_15_y_source_ram_renable <= 0;
        _mul_15_y_source_fifo_deq <= 0;
      end 
      _mul_15_y_idle <= _mul_15_y_idle;
      if(_mul_15_stream_oready) begin
        _mul_15_rshift_source_ram_renable <= 0;
        _mul_15_rshift_source_fifo_deq <= 0;
      end 
      _mul_15_rshift_idle <= _mul_15_rshift_idle;
      if(_mul_15_stream_oready) begin
        _mul_15_z_sink_wenable <= 0;
        _mul_15_z_sink_fifo_enq <= 0;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_1 <= _mul_15_stream_ivalid;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_2 <= __mul_15_stream_ivalid_1;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_3 <= __mul_15_stream_ivalid_2;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_4 <= __mul_15_stream_ivalid_3;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_5 <= __mul_15_stream_ivalid_4;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_6 <= __mul_15_stream_ivalid_5;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_7 <= __mul_15_stream_ivalid_6;
      end 
      if(_mul_15_stream_oready) begin
        __mul_15_stream_ivalid_8 <= __mul_15_stream_ivalid_7;
      end 
      if(_mul_15_stream_oready) begin
        _greaterthan_data_326 <= mul_15_rshift_data > 1'sd0;
      end 
      if(_mul_15_stream_oready) begin
        _minus_data_328 <= mul_15_rshift_data - 2'sd1;
      end 
      if(_mul_15_stream_oready) begin
        _greatereq_data_339 <= mul_15_x_data >= 1'sd0;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1735__variable_323 <= mul_15_x_data;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1738__variable_324 <= mul_15_y_data;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1741__variable_325 <= mul_15_rshift_data;
      end 
      if(_mul_15_stream_oready) begin
        _sll_data_330 <= 2'sd1 << _minus_data_328;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1732_greaterthan_326 <= _greaterthan_data_326;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1733_greatereq_339 <= _greatereq_data_339;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1736__delay_1735__variable_323 <= __delay_data_1735__variable_323;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1739__delay_1738__variable_324 <= __delay_data_1738__variable_324;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1742__delay_1741__variable_325 <= __delay_data_1741__variable_325;
      end 
      if(_mul_15_stream_oready) begin
        _cond_data_336 <= (__delay_data_1732_greaterthan_326)? _sll_data_330 : 1'sd0;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1734__delay_1733_greatereq_339 <= __delay_data_1733_greatereq_339;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1737__delay_1736__delay_1735__variable_323 <= __delay_data_1736__delay_1735__variable_323;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1740__delay_1739__delay_1738__variable_324 <= __delay_data_1739__delay_1738__variable_324;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1743__delay_1742__delay_1741__variable_325 <= __delay_data_1742__delay_1741__variable_325;
      end 
      if(_mul_15_stream_oready) begin
        __muladd_madd_odata_reg_342 <= __muladd_madd_odata_342;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1744__delay_1743__delay_1742____variable_325 <= __delay_data_1743__delay_1742__delay_1741__variable_325;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1745__delay_1744__delay_1743____variable_325 <= __delay_data_1744__delay_1743__delay_1742____variable_325;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1746__delay_1745__delay_1744____variable_325 <= __delay_data_1745__delay_1744__delay_1743____variable_325;
      end 
      if(_mul_15_stream_oready) begin
        __delay_data_1747__delay_1746__delay_1745____variable_325 <= __delay_data_1746__delay_1745__delay_1744____variable_325;
      end 
      if(_mul_15_stream_oready) begin
        _sra_data_343 <= __muladd_data_342 >>> __delay_data_1747__delay_1746__delay_1745____variable_325;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_323 <= _cond_data_1595;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_324 <= _cond_data_1433;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_325 <= __delay_data_2783__delay_2782_plus_1748;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_726 <= _mul_15_source_start;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_727 <= _tmp_726;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_728 <= _tmp_727;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_729 <= _mul_15_source_start;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_730 <= _tmp_729;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_731 <= _tmp_730;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_732 <= _tmp_731;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_733 <= _tmp_732;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_734 <= _tmp_733;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_735 <= _tmp_734;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_736 <= _tmp_735;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_737 <= _tmp_736;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_738 <= _tmp_737;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_739 <= _mul_15_source_stop;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_740 <= _tmp_739;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_741 <= _tmp_740;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_742 <= _tmp_741;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_743 <= _tmp_742;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_744 <= _tmp_743;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_745 <= _tmp_744;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_746 <= _tmp_745;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_747 <= _tmp_746;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_748 <= _tmp_747;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_749 <= _mul_15_source_busy;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_750 <= _tmp_749;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_751 <= _tmp_750;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_752 <= _tmp_751;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_753 <= _tmp_752;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_754 <= _tmp_753;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_755 <= _tmp_754;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_756 <= _tmp_755;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_757 <= _tmp_756;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_758 <= _tmp_757;
      end 
      if(_mul_15_stream_oready) begin
        _tmp_759 <= _mul_15_sink_busy;
      end 
      if(!_mul_15_sink_busy && _tmp_759) begin
        _mul_15_busy_reg <= 0;
      end 
      if(_mul_15_source_busy) begin
        _mul_15_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_15_fsm_1 = 1;
  localparam _mul_15_fsm_2 = 2;
  localparam _mul_15_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_15_fsm <= _mul_15_fsm_init;
      _mul_15_source_start <= 0;
      _mul_15_source_busy <= 0;
      _mul_15_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_15_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_15_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_15_stream_oready && _tmp_728) begin
        _mul_15_stream_ivalid <= 1;
      end 
      if(_mul_15_stream_oready && 1'd0) begin
        _mul_15_stream_ivalid <= 0;
      end 
      case(_mul_15_fsm)
        _mul_15_fsm_init: begin
          if(_mul_15_run_flag) begin
            _mul_15_source_start <= 1;
          end 
          if(_mul_15_run_flag) begin
            _mul_15_fsm <= _mul_15_fsm_1;
          end 
        end
        _mul_15_fsm_1: begin
          if(_mul_15_source_start && _mul_15_stream_oready) begin
            _mul_15_source_start <= 0;
            _mul_15_source_busy <= 1;
          end 
          if(_mul_15_source_start && _mul_15_stream_oready) begin
            _mul_15_fsm <= _mul_15_fsm_2;
          end 
        end
        _mul_15_fsm_2: begin
          if(_mul_15_stream_oready) begin
            _mul_15_fsm <= _mul_15_fsm_3;
          end 
        end
        _mul_15_fsm_3: begin
          if(_mul_15_stream_oready && 1'd0) begin
            _mul_15_source_busy <= 0;
          end 
          if(_mul_15_stream_oready && 1'd0 && _mul_15_run_flag) begin
            _mul_15_source_start <= 1;
          end 
          if(_mul_15_stream_oready && 1'd0) begin
            _mul_15_fsm <= _mul_15_fsm_init;
          end 
          if(_mul_15_stream_oready && 1'd0 && _mul_15_run_flag) begin
            _mul_15_fsm <= _mul_15_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_16_x_source_ram_renable <= 0;
      _mul_16_x_source_fifo_deq <= 0;
      _mul_16_x_idle <= 1;
      _mul_16_y_source_ram_renable <= 0;
      _mul_16_y_source_fifo_deq <= 0;
      _mul_16_y_idle <= 1;
      _mul_16_rshift_source_ram_renable <= 0;
      _mul_16_rshift_source_fifo_deq <= 0;
      _mul_16_rshift_idle <= 1;
      _mul_16_z_sink_wenable <= 0;
      _mul_16_z_sink_fifo_enq <= 0;
      __mul_16_stream_ivalid_1 <= 0;
      __mul_16_stream_ivalid_2 <= 0;
      __mul_16_stream_ivalid_3 <= 0;
      __mul_16_stream_ivalid_4 <= 0;
      __mul_16_stream_ivalid_5 <= 0;
      __mul_16_stream_ivalid_6 <= 0;
      __mul_16_stream_ivalid_7 <= 0;
      __mul_16_stream_ivalid_8 <= 0;
      _greaterthan_data_347 <= 0;
      _minus_data_349 <= 0;
      _greatereq_data_360 <= 0;
      __delay_data_1754__variable_344 <= 0;
      __delay_data_1757__variable_345 <= 0;
      __delay_data_1760__variable_346 <= 0;
      _sll_data_351 <= 0;
      __delay_data_1751_greaterthan_347 <= 0;
      __delay_data_1752_greatereq_360 <= 0;
      __delay_data_1755__delay_1754__variable_344 <= 0;
      __delay_data_1758__delay_1757__variable_345 <= 0;
      __delay_data_1761__delay_1760__variable_346 <= 0;
      _cond_data_357 <= 0;
      __delay_data_1753__delay_1752_greatereq_360 <= 0;
      __delay_data_1756__delay_1755__delay_1754__variable_344 <= 0;
      __delay_data_1759__delay_1758__delay_1757__variable_345 <= 0;
      __delay_data_1762__delay_1761__delay_1760__variable_346 <= 0;
      __muladd_madd_odata_reg_363 <= 0;
      __delay_data_1763__delay_1762__delay_1761____variable_346 <= 0;
      __delay_data_1764__delay_1763__delay_1762____variable_346 <= 0;
      __delay_data_1765__delay_1764__delay_1763____variable_346 <= 0;
      __delay_data_1766__delay_1765__delay_1764____variable_346 <= 0;
      _sra_data_364 <= 0;
      __variable_wdata_344 <= 0;
      __variable_wdata_345 <= 0;
      __variable_wdata_346 <= 0;
      _tmp_760 <= 0;
      _tmp_761 <= 0;
      _tmp_762 <= 0;
      _tmp_763 <= 0;
      _tmp_764 <= 0;
      _tmp_765 <= 0;
      _tmp_766 <= 0;
      _tmp_767 <= 0;
      _tmp_768 <= 0;
      _tmp_769 <= 0;
      _tmp_770 <= 0;
      _tmp_771 <= 0;
      _tmp_772 <= 0;
      _tmp_773 <= 0;
      _tmp_774 <= 0;
      _tmp_775 <= 0;
      _tmp_776 <= 0;
      _tmp_777 <= 0;
      _tmp_778 <= 0;
      _tmp_779 <= 0;
      _tmp_780 <= 0;
      _tmp_781 <= 0;
      _tmp_782 <= 0;
      _tmp_783 <= 0;
      _tmp_784 <= 0;
      _tmp_785 <= 0;
      _tmp_786 <= 0;
      _tmp_787 <= 0;
      _tmp_788 <= 0;
      _tmp_789 <= 0;
      _tmp_790 <= 0;
      _tmp_791 <= 0;
      _tmp_792 <= 0;
      _tmp_793 <= 0;
      _mul_16_busy_reg <= 0;
    end else begin
      if(_mul_16_stream_oready) begin
        _mul_16_x_source_ram_renable <= 0;
        _mul_16_x_source_fifo_deq <= 0;
      end 
      _mul_16_x_idle <= _mul_16_x_idle;
      if(_mul_16_stream_oready) begin
        _mul_16_y_source_ram_renable <= 0;
        _mul_16_y_source_fifo_deq <= 0;
      end 
      _mul_16_y_idle <= _mul_16_y_idle;
      if(_mul_16_stream_oready) begin
        _mul_16_rshift_source_ram_renable <= 0;
        _mul_16_rshift_source_fifo_deq <= 0;
      end 
      _mul_16_rshift_idle <= _mul_16_rshift_idle;
      if(_mul_16_stream_oready) begin
        _mul_16_z_sink_wenable <= 0;
        _mul_16_z_sink_fifo_enq <= 0;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_1 <= _mul_16_stream_ivalid;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_2 <= __mul_16_stream_ivalid_1;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_3 <= __mul_16_stream_ivalid_2;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_4 <= __mul_16_stream_ivalid_3;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_5 <= __mul_16_stream_ivalid_4;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_6 <= __mul_16_stream_ivalid_5;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_7 <= __mul_16_stream_ivalid_6;
      end 
      if(_mul_16_stream_oready) begin
        __mul_16_stream_ivalid_8 <= __mul_16_stream_ivalid_7;
      end 
      if(_mul_16_stream_oready) begin
        _greaterthan_data_347 <= mul_16_rshift_data > 1'sd0;
      end 
      if(_mul_16_stream_oready) begin
        _minus_data_349 <= mul_16_rshift_data - 2'sd1;
      end 
      if(_mul_16_stream_oready) begin
        _greatereq_data_360 <= mul_16_x_data >= 1'sd0;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1754__variable_344 <= mul_16_x_data;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1757__variable_345 <= mul_16_y_data;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1760__variable_346 <= mul_16_rshift_data;
      end 
      if(_mul_16_stream_oready) begin
        _sll_data_351 <= 2'sd1 << _minus_data_349;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1751_greaterthan_347 <= _greaterthan_data_347;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1752_greatereq_360 <= _greatereq_data_360;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1755__delay_1754__variable_344 <= __delay_data_1754__variable_344;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1758__delay_1757__variable_345 <= __delay_data_1757__variable_345;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1761__delay_1760__variable_346 <= __delay_data_1760__variable_346;
      end 
      if(_mul_16_stream_oready) begin
        _cond_data_357 <= (__delay_data_1751_greaterthan_347)? _sll_data_351 : 1'sd0;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1753__delay_1752_greatereq_360 <= __delay_data_1752_greatereq_360;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1756__delay_1755__delay_1754__variable_344 <= __delay_data_1755__delay_1754__variable_344;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1759__delay_1758__delay_1757__variable_345 <= __delay_data_1758__delay_1757__variable_345;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1762__delay_1761__delay_1760__variable_346 <= __delay_data_1761__delay_1760__variable_346;
      end 
      if(_mul_16_stream_oready) begin
        __muladd_madd_odata_reg_363 <= __muladd_madd_odata_363;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1763__delay_1762__delay_1761____variable_346 <= __delay_data_1762__delay_1761__delay_1760__variable_346;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1764__delay_1763__delay_1762____variable_346 <= __delay_data_1763__delay_1762__delay_1761____variable_346;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1765__delay_1764__delay_1763____variable_346 <= __delay_data_1764__delay_1763__delay_1762____variable_346;
      end 
      if(_mul_16_stream_oready) begin
        __delay_data_1766__delay_1765__delay_1764____variable_346 <= __delay_data_1765__delay_1764__delay_1763____variable_346;
      end 
      if(_mul_16_stream_oready) begin
        _sra_data_364 <= __muladd_data_363 >>> __delay_data_1766__delay_1765__delay_1764____variable_346;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_344 <= _cond_data_1597;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_345 <= _cond_data_1435;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_346 <= __delay_data_2800__delay_2799_plus_1767;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_760 <= _mul_16_source_start;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_761 <= _tmp_760;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_762 <= _tmp_761;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_763 <= _mul_16_source_start;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_764 <= _tmp_763;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_765 <= _tmp_764;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_766 <= _tmp_765;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_767 <= _tmp_766;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_768 <= _tmp_767;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_769 <= _tmp_768;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_770 <= _tmp_769;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_771 <= _tmp_770;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_772 <= _tmp_771;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_773 <= _mul_16_source_stop;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_774 <= _tmp_773;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_775 <= _tmp_774;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_776 <= _tmp_775;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_777 <= _tmp_776;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_778 <= _tmp_777;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_779 <= _tmp_778;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_780 <= _tmp_779;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_781 <= _tmp_780;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_782 <= _tmp_781;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_783 <= _mul_16_source_busy;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_784 <= _tmp_783;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_785 <= _tmp_784;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_786 <= _tmp_785;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_787 <= _tmp_786;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_788 <= _tmp_787;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_789 <= _tmp_788;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_790 <= _tmp_789;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_791 <= _tmp_790;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_792 <= _tmp_791;
      end 
      if(_mul_16_stream_oready) begin
        _tmp_793 <= _mul_16_sink_busy;
      end 
      if(!_mul_16_sink_busy && _tmp_793) begin
        _mul_16_busy_reg <= 0;
      end 
      if(_mul_16_source_busy) begin
        _mul_16_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_16_fsm_1 = 1;
  localparam _mul_16_fsm_2 = 2;
  localparam _mul_16_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_16_fsm <= _mul_16_fsm_init;
      _mul_16_source_start <= 0;
      _mul_16_source_busy <= 0;
      _mul_16_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_16_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_16_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_16_stream_oready && _tmp_762) begin
        _mul_16_stream_ivalid <= 1;
      end 
      if(_mul_16_stream_oready && 1'd0) begin
        _mul_16_stream_ivalid <= 0;
      end 
      case(_mul_16_fsm)
        _mul_16_fsm_init: begin
          if(_mul_16_run_flag) begin
            _mul_16_source_start <= 1;
          end 
          if(_mul_16_run_flag) begin
            _mul_16_fsm <= _mul_16_fsm_1;
          end 
        end
        _mul_16_fsm_1: begin
          if(_mul_16_source_start && _mul_16_stream_oready) begin
            _mul_16_source_start <= 0;
            _mul_16_source_busy <= 1;
          end 
          if(_mul_16_source_start && _mul_16_stream_oready) begin
            _mul_16_fsm <= _mul_16_fsm_2;
          end 
        end
        _mul_16_fsm_2: begin
          if(_mul_16_stream_oready) begin
            _mul_16_fsm <= _mul_16_fsm_3;
          end 
        end
        _mul_16_fsm_3: begin
          if(_mul_16_stream_oready && 1'd0) begin
            _mul_16_source_busy <= 0;
          end 
          if(_mul_16_stream_oready && 1'd0 && _mul_16_run_flag) begin
            _mul_16_source_start <= 1;
          end 
          if(_mul_16_stream_oready && 1'd0) begin
            _mul_16_fsm <= _mul_16_fsm_init;
          end 
          if(_mul_16_stream_oready && 1'd0 && _mul_16_run_flag) begin
            _mul_16_fsm <= _mul_16_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_17_x_source_ram_renable <= 0;
      _mul_17_x_source_fifo_deq <= 0;
      _mul_17_x_idle <= 1;
      _mul_17_y_source_ram_renable <= 0;
      _mul_17_y_source_fifo_deq <= 0;
      _mul_17_y_idle <= 1;
      _mul_17_rshift_source_ram_renable <= 0;
      _mul_17_rshift_source_fifo_deq <= 0;
      _mul_17_rshift_idle <= 1;
      _mul_17_z_sink_wenable <= 0;
      _mul_17_z_sink_fifo_enq <= 0;
      __mul_17_stream_ivalid_1 <= 0;
      __mul_17_stream_ivalid_2 <= 0;
      __mul_17_stream_ivalid_3 <= 0;
      __mul_17_stream_ivalid_4 <= 0;
      __mul_17_stream_ivalid_5 <= 0;
      __mul_17_stream_ivalid_6 <= 0;
      __mul_17_stream_ivalid_7 <= 0;
      __mul_17_stream_ivalid_8 <= 0;
      _greaterthan_data_368 <= 0;
      _minus_data_370 <= 0;
      _greatereq_data_381 <= 0;
      __delay_data_1791__variable_365 <= 0;
      __delay_data_1794__variable_366 <= 0;
      __delay_data_1797__variable_367 <= 0;
      _sll_data_372 <= 0;
      __delay_data_1788_greaterthan_368 <= 0;
      __delay_data_1789_greatereq_381 <= 0;
      __delay_data_1792__delay_1791__variable_365 <= 0;
      __delay_data_1795__delay_1794__variable_366 <= 0;
      __delay_data_1798__delay_1797__variable_367 <= 0;
      _cond_data_378 <= 0;
      __delay_data_1790__delay_1789_greatereq_381 <= 0;
      __delay_data_1793__delay_1792__delay_1791__variable_365 <= 0;
      __delay_data_1796__delay_1795__delay_1794__variable_366 <= 0;
      __delay_data_1799__delay_1798__delay_1797__variable_367 <= 0;
      __muladd_madd_odata_reg_384 <= 0;
      __delay_data_1800__delay_1799__delay_1798____variable_367 <= 0;
      __delay_data_1801__delay_1800__delay_1799____variable_367 <= 0;
      __delay_data_1802__delay_1801__delay_1800____variable_367 <= 0;
      __delay_data_1803__delay_1802__delay_1801____variable_367 <= 0;
      _sra_data_385 <= 0;
      __variable_wdata_365 <= 0;
      __variable_wdata_366 <= 0;
      __variable_wdata_367 <= 0;
      _tmp_794 <= 0;
      _tmp_795 <= 0;
      _tmp_796 <= 0;
      _tmp_797 <= 0;
      _tmp_798 <= 0;
      _tmp_799 <= 0;
      _tmp_800 <= 0;
      _tmp_801 <= 0;
      _tmp_802 <= 0;
      _tmp_803 <= 0;
      _tmp_804 <= 0;
      _tmp_805 <= 0;
      _tmp_806 <= 0;
      _tmp_807 <= 0;
      _tmp_808 <= 0;
      _tmp_809 <= 0;
      _tmp_810 <= 0;
      _tmp_811 <= 0;
      _tmp_812 <= 0;
      _tmp_813 <= 0;
      _tmp_814 <= 0;
      _tmp_815 <= 0;
      _tmp_816 <= 0;
      _tmp_817 <= 0;
      _tmp_818 <= 0;
      _tmp_819 <= 0;
      _tmp_820 <= 0;
      _tmp_821 <= 0;
      _tmp_822 <= 0;
      _tmp_823 <= 0;
      _tmp_824 <= 0;
      _tmp_825 <= 0;
      _tmp_826 <= 0;
      _tmp_827 <= 0;
      _mul_17_busy_reg <= 0;
    end else begin
      if(_mul_17_stream_oready) begin
        _mul_17_x_source_ram_renable <= 0;
        _mul_17_x_source_fifo_deq <= 0;
      end 
      _mul_17_x_idle <= _mul_17_x_idle;
      if(_mul_17_stream_oready) begin
        _mul_17_y_source_ram_renable <= 0;
        _mul_17_y_source_fifo_deq <= 0;
      end 
      _mul_17_y_idle <= _mul_17_y_idle;
      if(_mul_17_stream_oready) begin
        _mul_17_rshift_source_ram_renable <= 0;
        _mul_17_rshift_source_fifo_deq <= 0;
      end 
      _mul_17_rshift_idle <= _mul_17_rshift_idle;
      if(_mul_17_stream_oready) begin
        _mul_17_z_sink_wenable <= 0;
        _mul_17_z_sink_fifo_enq <= 0;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_1 <= _mul_17_stream_ivalid;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_2 <= __mul_17_stream_ivalid_1;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_3 <= __mul_17_stream_ivalid_2;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_4 <= __mul_17_stream_ivalid_3;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_5 <= __mul_17_stream_ivalid_4;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_6 <= __mul_17_stream_ivalid_5;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_7 <= __mul_17_stream_ivalid_6;
      end 
      if(_mul_17_stream_oready) begin
        __mul_17_stream_ivalid_8 <= __mul_17_stream_ivalid_7;
      end 
      if(_mul_17_stream_oready) begin
        _greaterthan_data_368 <= mul_17_rshift_data > 1'sd0;
      end 
      if(_mul_17_stream_oready) begin
        _minus_data_370 <= mul_17_rshift_data - 2'sd1;
      end 
      if(_mul_17_stream_oready) begin
        _greatereq_data_381 <= mul_17_x_data >= 1'sd0;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1791__variable_365 <= mul_17_x_data;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1794__variable_366 <= mul_17_y_data;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1797__variable_367 <= mul_17_rshift_data;
      end 
      if(_mul_17_stream_oready) begin
        _sll_data_372 <= 2'sd1 << _minus_data_370;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1788_greaterthan_368 <= _greaterthan_data_368;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1789_greatereq_381 <= _greatereq_data_381;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1792__delay_1791__variable_365 <= __delay_data_1791__variable_365;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1795__delay_1794__variable_366 <= __delay_data_1794__variable_366;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1798__delay_1797__variable_367 <= __delay_data_1797__variable_367;
      end 
      if(_mul_17_stream_oready) begin
        _cond_data_378 <= (__delay_data_1788_greaterthan_368)? _sll_data_372 : 1'sd0;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1790__delay_1789_greatereq_381 <= __delay_data_1789_greatereq_381;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1793__delay_1792__delay_1791__variable_365 <= __delay_data_1792__delay_1791__variable_365;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1796__delay_1795__delay_1794__variable_366 <= __delay_data_1795__delay_1794__variable_366;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1799__delay_1798__delay_1797__variable_367 <= __delay_data_1798__delay_1797__variable_367;
      end 
      if(_mul_17_stream_oready) begin
        __muladd_madd_odata_reg_384 <= __muladd_madd_odata_384;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1800__delay_1799__delay_1798____variable_367 <= __delay_data_1799__delay_1798__delay_1797__variable_367;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1801__delay_1800__delay_1799____variable_367 <= __delay_data_1800__delay_1799__delay_1798____variable_367;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1802__delay_1801__delay_1800____variable_367 <= __delay_data_1801__delay_1800__delay_1799____variable_367;
      end 
      if(_mul_17_stream_oready) begin
        __delay_data_1803__delay_1802__delay_1801____variable_367 <= __delay_data_1802__delay_1801__delay_1800____variable_367;
      end 
      if(_mul_17_stream_oready) begin
        _sra_data_385 <= __muladd_data_384 >>> __delay_data_1803__delay_1802__delay_1801____variable_367;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_365 <= _cond_data_1770;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_366 <= _cond_data_1437;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_367 <= __delay_data_2671__delay_2670_plus_1804;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_794 <= _mul_17_source_start;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_795 <= _tmp_794;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_796 <= _tmp_795;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_797 <= _mul_17_source_start;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_798 <= _tmp_797;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_799 <= _tmp_798;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_800 <= _tmp_799;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_801 <= _tmp_800;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_802 <= _tmp_801;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_803 <= _tmp_802;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_804 <= _tmp_803;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_805 <= _tmp_804;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_806 <= _tmp_805;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_807 <= _mul_17_source_stop;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_808 <= _tmp_807;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_809 <= _tmp_808;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_810 <= _tmp_809;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_811 <= _tmp_810;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_812 <= _tmp_811;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_813 <= _tmp_812;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_814 <= _tmp_813;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_815 <= _tmp_814;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_816 <= _tmp_815;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_817 <= _mul_17_source_busy;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_818 <= _tmp_817;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_819 <= _tmp_818;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_820 <= _tmp_819;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_821 <= _tmp_820;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_822 <= _tmp_821;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_823 <= _tmp_822;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_824 <= _tmp_823;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_825 <= _tmp_824;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_826 <= _tmp_825;
      end 
      if(_mul_17_stream_oready) begin
        _tmp_827 <= _mul_17_sink_busy;
      end 
      if(!_mul_17_sink_busy && _tmp_827) begin
        _mul_17_busy_reg <= 0;
      end 
      if(_mul_17_source_busy) begin
        _mul_17_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_17_fsm_1 = 1;
  localparam _mul_17_fsm_2 = 2;
  localparam _mul_17_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_17_fsm <= _mul_17_fsm_init;
      _mul_17_source_start <= 0;
      _mul_17_source_busy <= 0;
      _mul_17_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_17_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_17_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_17_stream_oready && _tmp_796) begin
        _mul_17_stream_ivalid <= 1;
      end 
      if(_mul_17_stream_oready && 1'd0) begin
        _mul_17_stream_ivalid <= 0;
      end 
      case(_mul_17_fsm)
        _mul_17_fsm_init: begin
          if(_mul_17_run_flag) begin
            _mul_17_source_start <= 1;
          end 
          if(_mul_17_run_flag) begin
            _mul_17_fsm <= _mul_17_fsm_1;
          end 
        end
        _mul_17_fsm_1: begin
          if(_mul_17_source_start && _mul_17_stream_oready) begin
            _mul_17_source_start <= 0;
            _mul_17_source_busy <= 1;
          end 
          if(_mul_17_source_start && _mul_17_stream_oready) begin
            _mul_17_fsm <= _mul_17_fsm_2;
          end 
        end
        _mul_17_fsm_2: begin
          if(_mul_17_stream_oready) begin
            _mul_17_fsm <= _mul_17_fsm_3;
          end 
        end
        _mul_17_fsm_3: begin
          if(_mul_17_stream_oready && 1'd0) begin
            _mul_17_source_busy <= 0;
          end 
          if(_mul_17_stream_oready && 1'd0 && _mul_17_run_flag) begin
            _mul_17_source_start <= 1;
          end 
          if(_mul_17_stream_oready && 1'd0) begin
            _mul_17_fsm <= _mul_17_fsm_init;
          end 
          if(_mul_17_stream_oready && 1'd0 && _mul_17_run_flag) begin
            _mul_17_fsm <= _mul_17_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_18_x_source_ram_renable <= 0;
      _mul_18_x_source_fifo_deq <= 0;
      _mul_18_x_idle <= 1;
      _mul_18_y_source_ram_renable <= 0;
      _mul_18_y_source_fifo_deq <= 0;
      _mul_18_y_idle <= 1;
      _mul_18_rshift_source_ram_renable <= 0;
      _mul_18_rshift_source_fifo_deq <= 0;
      _mul_18_rshift_idle <= 1;
      _mul_18_z_sink_wenable <= 0;
      _mul_18_z_sink_fifo_enq <= 0;
      __mul_18_stream_ivalid_1 <= 0;
      __mul_18_stream_ivalid_2 <= 0;
      __mul_18_stream_ivalid_3 <= 0;
      __mul_18_stream_ivalid_4 <= 0;
      __mul_18_stream_ivalid_5 <= 0;
      __mul_18_stream_ivalid_6 <= 0;
      __mul_18_stream_ivalid_7 <= 0;
      __mul_18_stream_ivalid_8 <= 0;
      _greaterthan_data_389 <= 0;
      _minus_data_391 <= 0;
      _greatereq_data_402 <= 0;
      __delay_data_1810__variable_386 <= 0;
      __delay_data_1813__variable_387 <= 0;
      __delay_data_1816__variable_388 <= 0;
      _sll_data_393 <= 0;
      __delay_data_1807_greaterthan_389 <= 0;
      __delay_data_1808_greatereq_402 <= 0;
      __delay_data_1811__delay_1810__variable_386 <= 0;
      __delay_data_1814__delay_1813__variable_387 <= 0;
      __delay_data_1817__delay_1816__variable_388 <= 0;
      _cond_data_399 <= 0;
      __delay_data_1809__delay_1808_greatereq_402 <= 0;
      __delay_data_1812__delay_1811__delay_1810__variable_386 <= 0;
      __delay_data_1815__delay_1814__delay_1813__variable_387 <= 0;
      __delay_data_1818__delay_1817__delay_1816__variable_388 <= 0;
      __muladd_madd_odata_reg_405 <= 0;
      __delay_data_1819__delay_1818__delay_1817____variable_388 <= 0;
      __delay_data_1820__delay_1819__delay_1818____variable_388 <= 0;
      __delay_data_1821__delay_1820__delay_1819____variable_388 <= 0;
      __delay_data_1822__delay_1821__delay_1820____variable_388 <= 0;
      _sra_data_406 <= 0;
      __variable_wdata_386 <= 0;
      __variable_wdata_387 <= 0;
      __variable_wdata_388 <= 0;
      _tmp_828 <= 0;
      _tmp_829 <= 0;
      _tmp_830 <= 0;
      _tmp_831 <= 0;
      _tmp_832 <= 0;
      _tmp_833 <= 0;
      _tmp_834 <= 0;
      _tmp_835 <= 0;
      _tmp_836 <= 0;
      _tmp_837 <= 0;
      _tmp_838 <= 0;
      _tmp_839 <= 0;
      _tmp_840 <= 0;
      _tmp_841 <= 0;
      _tmp_842 <= 0;
      _tmp_843 <= 0;
      _tmp_844 <= 0;
      _tmp_845 <= 0;
      _tmp_846 <= 0;
      _tmp_847 <= 0;
      _tmp_848 <= 0;
      _tmp_849 <= 0;
      _tmp_850 <= 0;
      _tmp_851 <= 0;
      _tmp_852 <= 0;
      _tmp_853 <= 0;
      _tmp_854 <= 0;
      _tmp_855 <= 0;
      _tmp_856 <= 0;
      _tmp_857 <= 0;
      _tmp_858 <= 0;
      _tmp_859 <= 0;
      _tmp_860 <= 0;
      _tmp_861 <= 0;
      _mul_18_busy_reg <= 0;
    end else begin
      if(_mul_18_stream_oready) begin
        _mul_18_x_source_ram_renable <= 0;
        _mul_18_x_source_fifo_deq <= 0;
      end 
      _mul_18_x_idle <= _mul_18_x_idle;
      if(_mul_18_stream_oready) begin
        _mul_18_y_source_ram_renable <= 0;
        _mul_18_y_source_fifo_deq <= 0;
      end 
      _mul_18_y_idle <= _mul_18_y_idle;
      if(_mul_18_stream_oready) begin
        _mul_18_rshift_source_ram_renable <= 0;
        _mul_18_rshift_source_fifo_deq <= 0;
      end 
      _mul_18_rshift_idle <= _mul_18_rshift_idle;
      if(_mul_18_stream_oready) begin
        _mul_18_z_sink_wenable <= 0;
        _mul_18_z_sink_fifo_enq <= 0;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_1 <= _mul_18_stream_ivalid;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_2 <= __mul_18_stream_ivalid_1;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_3 <= __mul_18_stream_ivalid_2;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_4 <= __mul_18_stream_ivalid_3;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_5 <= __mul_18_stream_ivalid_4;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_6 <= __mul_18_stream_ivalid_5;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_7 <= __mul_18_stream_ivalid_6;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_8 <= __mul_18_stream_ivalid_7;
      end 
      if(_mul_18_stream_oready) begin
        _greaterthan_data_389 <= mul_18_rshift_data > 1'sd0;
      end 
      if(_mul_18_stream_oready) begin
        _minus_data_391 <= mul_18_rshift_data - 2'sd1;
      end 
      if(_mul_18_stream_oready) begin
        _greatereq_data_402 <= mul_18_x_data >= 1'sd0;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1810__variable_386 <= mul_18_x_data;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1813__variable_387 <= mul_18_y_data;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1816__variable_388 <= mul_18_rshift_data;
      end 
      if(_mul_18_stream_oready) begin
        _sll_data_393 <= 2'sd1 << _minus_data_391;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1807_greaterthan_389 <= _greaterthan_data_389;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1808_greatereq_402 <= _greatereq_data_402;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1811__delay_1810__variable_386 <= __delay_data_1810__variable_386;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1814__delay_1813__variable_387 <= __delay_data_1813__variable_387;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1817__delay_1816__variable_388 <= __delay_data_1816__variable_388;
      end 
      if(_mul_18_stream_oready) begin
        _cond_data_399 <= (__delay_data_1807_greaterthan_389)? _sll_data_393 : 1'sd0;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1809__delay_1808_greatereq_402 <= __delay_data_1808_greatereq_402;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1812__delay_1811__delay_1810__variable_386 <= __delay_data_1811__delay_1810__variable_386;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1815__delay_1814__delay_1813__variable_387 <= __delay_data_1814__delay_1813__variable_387;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1818__delay_1817__delay_1816__variable_388 <= __delay_data_1817__delay_1816__variable_388;
      end 
      if(_mul_18_stream_oready) begin
        __muladd_madd_odata_reg_405 <= __muladd_madd_odata_405;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1819__delay_1818__delay_1817____variable_388 <= __delay_data_1818__delay_1817__delay_1816__variable_388;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1820__delay_1819__delay_1818____variable_388 <= __delay_data_1819__delay_1818__delay_1817____variable_388;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1821__delay_1820__delay_1819____variable_388 <= __delay_data_1820__delay_1819__delay_1818____variable_388;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1822__delay_1821__delay_1820____variable_388 <= __delay_data_1821__delay_1820__delay_1819____variable_388;
      end 
      if(_mul_18_stream_oready) begin
        _sra_data_406 <= __muladd_data_405 >>> __delay_data_1822__delay_1821__delay_1820____variable_388;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_386 <= _cond_data_1772;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_387 <= _cond_data_1439;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_388 <= __delay_data_2688__delay_2687_plus_1823;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_828 <= _mul_18_source_start;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_829 <= _tmp_828;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_830 <= _tmp_829;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_831 <= _mul_18_source_start;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_832 <= _tmp_831;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_833 <= _tmp_832;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_834 <= _tmp_833;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_835 <= _tmp_834;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_836 <= _tmp_835;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_837 <= _tmp_836;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_838 <= _tmp_837;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_839 <= _tmp_838;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_840 <= _tmp_839;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_841 <= _mul_18_source_stop;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_842 <= _tmp_841;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_843 <= _tmp_842;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_844 <= _tmp_843;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_845 <= _tmp_844;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_846 <= _tmp_845;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_847 <= _tmp_846;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_848 <= _tmp_847;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_849 <= _tmp_848;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_850 <= _tmp_849;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_851 <= _mul_18_source_busy;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_852 <= _tmp_851;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_853 <= _tmp_852;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_854 <= _tmp_853;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_855 <= _tmp_854;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_856 <= _tmp_855;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_857 <= _tmp_856;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_858 <= _tmp_857;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_859 <= _tmp_858;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_860 <= _tmp_859;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_861 <= _mul_18_sink_busy;
      end 
      if(!_mul_18_sink_busy && _tmp_861) begin
        _mul_18_busy_reg <= 0;
      end 
      if(_mul_18_source_busy) begin
        _mul_18_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_18_fsm_1 = 1;
  localparam _mul_18_fsm_2 = 2;
  localparam _mul_18_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_18_fsm <= _mul_18_fsm_init;
      _mul_18_source_start <= 0;
      _mul_18_source_busy <= 0;
      _mul_18_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_18_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_18_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_18_stream_oready && _tmp_830) begin
        _mul_18_stream_ivalid <= 1;
      end 
      if(_mul_18_stream_oready && 1'd0) begin
        _mul_18_stream_ivalid <= 0;
      end 
      case(_mul_18_fsm)
        _mul_18_fsm_init: begin
          if(_mul_18_run_flag) begin
            _mul_18_source_start <= 1;
          end 
          if(_mul_18_run_flag) begin
            _mul_18_fsm <= _mul_18_fsm_1;
          end 
        end
        _mul_18_fsm_1: begin
          if(_mul_18_source_start && _mul_18_stream_oready) begin
            _mul_18_source_start <= 0;
            _mul_18_source_busy <= 1;
          end 
          if(_mul_18_source_start && _mul_18_stream_oready) begin
            _mul_18_fsm <= _mul_18_fsm_2;
          end 
        end
        _mul_18_fsm_2: begin
          if(_mul_18_stream_oready) begin
            _mul_18_fsm <= _mul_18_fsm_3;
          end 
        end
        _mul_18_fsm_3: begin
          if(_mul_18_stream_oready && 1'd0) begin
            _mul_18_source_busy <= 0;
          end 
          if(_mul_18_stream_oready && 1'd0 && _mul_18_run_flag) begin
            _mul_18_source_start <= 1;
          end 
          if(_mul_18_stream_oready && 1'd0) begin
            _mul_18_fsm <= _mul_18_fsm_init;
          end 
          if(_mul_18_stream_oready && 1'd0 && _mul_18_run_flag) begin
            _mul_18_fsm <= _mul_18_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_19_x_source_ram_renable <= 0;
      _mul_19_x_source_fifo_deq <= 0;
      _mul_19_x_idle <= 1;
      _mul_19_y_source_ram_renable <= 0;
      _mul_19_y_source_fifo_deq <= 0;
      _mul_19_y_idle <= 1;
      _mul_19_rshift_source_ram_renable <= 0;
      _mul_19_rshift_source_fifo_deq <= 0;
      _mul_19_rshift_idle <= 1;
      _mul_19_z_sink_wenable <= 0;
      _mul_19_z_sink_fifo_enq <= 0;
      __mul_19_stream_ivalid_1 <= 0;
      __mul_19_stream_ivalid_2 <= 0;
      __mul_19_stream_ivalid_3 <= 0;
      __mul_19_stream_ivalid_4 <= 0;
      __mul_19_stream_ivalid_5 <= 0;
      __mul_19_stream_ivalid_6 <= 0;
      __mul_19_stream_ivalid_7 <= 0;
      __mul_19_stream_ivalid_8 <= 0;
      _greaterthan_data_410 <= 0;
      _minus_data_412 <= 0;
      _greatereq_data_423 <= 0;
      __delay_data_1829__variable_407 <= 0;
      __delay_data_1832__variable_408 <= 0;
      __delay_data_1835__variable_409 <= 0;
      _sll_data_414 <= 0;
      __delay_data_1826_greaterthan_410 <= 0;
      __delay_data_1827_greatereq_423 <= 0;
      __delay_data_1830__delay_1829__variable_407 <= 0;
      __delay_data_1833__delay_1832__variable_408 <= 0;
      __delay_data_1836__delay_1835__variable_409 <= 0;
      _cond_data_420 <= 0;
      __delay_data_1828__delay_1827_greatereq_423 <= 0;
      __delay_data_1831__delay_1830__delay_1829__variable_407 <= 0;
      __delay_data_1834__delay_1833__delay_1832__variable_408 <= 0;
      __delay_data_1837__delay_1836__delay_1835__variable_409 <= 0;
      __muladd_madd_odata_reg_426 <= 0;
      __delay_data_1838__delay_1837__delay_1836____variable_409 <= 0;
      __delay_data_1839__delay_1838__delay_1837____variable_409 <= 0;
      __delay_data_1840__delay_1839__delay_1838____variable_409 <= 0;
      __delay_data_1841__delay_1840__delay_1839____variable_409 <= 0;
      _sra_data_427 <= 0;
      __variable_wdata_407 <= 0;
      __variable_wdata_408 <= 0;
      __variable_wdata_409 <= 0;
      _tmp_862 <= 0;
      _tmp_863 <= 0;
      _tmp_864 <= 0;
      _tmp_865 <= 0;
      _tmp_866 <= 0;
      _tmp_867 <= 0;
      _tmp_868 <= 0;
      _tmp_869 <= 0;
      _tmp_870 <= 0;
      _tmp_871 <= 0;
      _tmp_872 <= 0;
      _tmp_873 <= 0;
      _tmp_874 <= 0;
      _tmp_875 <= 0;
      _tmp_876 <= 0;
      _tmp_877 <= 0;
      _tmp_878 <= 0;
      _tmp_879 <= 0;
      _tmp_880 <= 0;
      _tmp_881 <= 0;
      _tmp_882 <= 0;
      _tmp_883 <= 0;
      _tmp_884 <= 0;
      _tmp_885 <= 0;
      _tmp_886 <= 0;
      _tmp_887 <= 0;
      _tmp_888 <= 0;
      _tmp_889 <= 0;
      _tmp_890 <= 0;
      _tmp_891 <= 0;
      _tmp_892 <= 0;
      _tmp_893 <= 0;
      _tmp_894 <= 0;
      _tmp_895 <= 0;
      _mul_19_busy_reg <= 0;
    end else begin
      if(_mul_19_stream_oready) begin
        _mul_19_x_source_ram_renable <= 0;
        _mul_19_x_source_fifo_deq <= 0;
      end 
      _mul_19_x_idle <= _mul_19_x_idle;
      if(_mul_19_stream_oready) begin
        _mul_19_y_source_ram_renable <= 0;
        _mul_19_y_source_fifo_deq <= 0;
      end 
      _mul_19_y_idle <= _mul_19_y_idle;
      if(_mul_19_stream_oready) begin
        _mul_19_rshift_source_ram_renable <= 0;
        _mul_19_rshift_source_fifo_deq <= 0;
      end 
      _mul_19_rshift_idle <= _mul_19_rshift_idle;
      if(_mul_19_stream_oready) begin
        _mul_19_z_sink_wenable <= 0;
        _mul_19_z_sink_fifo_enq <= 0;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_1 <= _mul_19_stream_ivalid;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_2 <= __mul_19_stream_ivalid_1;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_3 <= __mul_19_stream_ivalid_2;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_4 <= __mul_19_stream_ivalid_3;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_5 <= __mul_19_stream_ivalid_4;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_6 <= __mul_19_stream_ivalid_5;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_7 <= __mul_19_stream_ivalid_6;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_8 <= __mul_19_stream_ivalid_7;
      end 
      if(_mul_19_stream_oready) begin
        _greaterthan_data_410 <= mul_19_rshift_data > 1'sd0;
      end 
      if(_mul_19_stream_oready) begin
        _minus_data_412 <= mul_19_rshift_data - 2'sd1;
      end 
      if(_mul_19_stream_oready) begin
        _greatereq_data_423 <= mul_19_x_data >= 1'sd0;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1829__variable_407 <= mul_19_x_data;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1832__variable_408 <= mul_19_y_data;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1835__variable_409 <= mul_19_rshift_data;
      end 
      if(_mul_19_stream_oready) begin
        _sll_data_414 <= 2'sd1 << _minus_data_412;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1826_greaterthan_410 <= _greaterthan_data_410;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1827_greatereq_423 <= _greatereq_data_423;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1830__delay_1829__variable_407 <= __delay_data_1829__variable_407;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1833__delay_1832__variable_408 <= __delay_data_1832__variable_408;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1836__delay_1835__variable_409 <= __delay_data_1835__variable_409;
      end 
      if(_mul_19_stream_oready) begin
        _cond_data_420 <= (__delay_data_1826_greaterthan_410)? _sll_data_414 : 1'sd0;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1828__delay_1827_greatereq_423 <= __delay_data_1827_greatereq_423;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1831__delay_1830__delay_1829__variable_407 <= __delay_data_1830__delay_1829__variable_407;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1834__delay_1833__delay_1832__variable_408 <= __delay_data_1833__delay_1832__variable_408;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1837__delay_1836__delay_1835__variable_409 <= __delay_data_1836__delay_1835__variable_409;
      end 
      if(_mul_19_stream_oready) begin
        __muladd_madd_odata_reg_426 <= __muladd_madd_odata_426;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1838__delay_1837__delay_1836____variable_409 <= __delay_data_1837__delay_1836__delay_1835__variable_409;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1839__delay_1838__delay_1837____variable_409 <= __delay_data_1838__delay_1837__delay_1836____variable_409;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1840__delay_1839__delay_1838____variable_409 <= __delay_data_1839__delay_1838__delay_1837____variable_409;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1841__delay_1840__delay_1839____variable_409 <= __delay_data_1840__delay_1839__delay_1838____variable_409;
      end 
      if(_mul_19_stream_oready) begin
        _sra_data_427 <= __muladd_data_426 >>> __delay_data_1841__delay_1840__delay_1839____variable_409;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_407 <= _cond_data_1774;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_408 <= _cond_data_1441;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_409 <= __delay_data_2705__delay_2704_plus_1842;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_862 <= _mul_19_source_start;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_863 <= _tmp_862;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_864 <= _tmp_863;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_865 <= _mul_19_source_start;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_866 <= _tmp_865;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_867 <= _tmp_866;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_868 <= _tmp_867;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_869 <= _tmp_868;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_870 <= _tmp_869;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_871 <= _tmp_870;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_872 <= _tmp_871;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_873 <= _tmp_872;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_874 <= _tmp_873;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_875 <= _mul_19_source_stop;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_876 <= _tmp_875;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_877 <= _tmp_876;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_878 <= _tmp_877;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_879 <= _tmp_878;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_880 <= _tmp_879;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_881 <= _tmp_880;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_882 <= _tmp_881;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_883 <= _tmp_882;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_884 <= _tmp_883;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_885 <= _mul_19_source_busy;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_886 <= _tmp_885;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_887 <= _tmp_886;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_888 <= _tmp_887;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_889 <= _tmp_888;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_890 <= _tmp_889;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_891 <= _tmp_890;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_892 <= _tmp_891;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_893 <= _tmp_892;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_894 <= _tmp_893;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_895 <= _mul_19_sink_busy;
      end 
      if(!_mul_19_sink_busy && _tmp_895) begin
        _mul_19_busy_reg <= 0;
      end 
      if(_mul_19_source_busy) begin
        _mul_19_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_19_fsm_1 = 1;
  localparam _mul_19_fsm_2 = 2;
  localparam _mul_19_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_19_fsm <= _mul_19_fsm_init;
      _mul_19_source_start <= 0;
      _mul_19_source_busy <= 0;
      _mul_19_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_19_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_19_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_19_stream_oready && _tmp_864) begin
        _mul_19_stream_ivalid <= 1;
      end 
      if(_mul_19_stream_oready && 1'd0) begin
        _mul_19_stream_ivalid <= 0;
      end 
      case(_mul_19_fsm)
        _mul_19_fsm_init: begin
          if(_mul_19_run_flag) begin
            _mul_19_source_start <= 1;
          end 
          if(_mul_19_run_flag) begin
            _mul_19_fsm <= _mul_19_fsm_1;
          end 
        end
        _mul_19_fsm_1: begin
          if(_mul_19_source_start && _mul_19_stream_oready) begin
            _mul_19_source_start <= 0;
            _mul_19_source_busy <= 1;
          end 
          if(_mul_19_source_start && _mul_19_stream_oready) begin
            _mul_19_fsm <= _mul_19_fsm_2;
          end 
        end
        _mul_19_fsm_2: begin
          if(_mul_19_stream_oready) begin
            _mul_19_fsm <= _mul_19_fsm_3;
          end 
        end
        _mul_19_fsm_3: begin
          if(_mul_19_stream_oready && 1'd0) begin
            _mul_19_source_busy <= 0;
          end 
          if(_mul_19_stream_oready && 1'd0 && _mul_19_run_flag) begin
            _mul_19_source_start <= 1;
          end 
          if(_mul_19_stream_oready && 1'd0) begin
            _mul_19_fsm <= _mul_19_fsm_init;
          end 
          if(_mul_19_stream_oready && 1'd0 && _mul_19_run_flag) begin
            _mul_19_fsm <= _mul_19_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_20_x_source_ram_renable <= 0;
      _mul_20_x_source_fifo_deq <= 0;
      _mul_20_x_idle <= 1;
      _mul_20_y_source_ram_renable <= 0;
      _mul_20_y_source_fifo_deq <= 0;
      _mul_20_y_idle <= 1;
      _mul_20_rshift_source_ram_renable <= 0;
      _mul_20_rshift_source_fifo_deq <= 0;
      _mul_20_rshift_idle <= 1;
      _mul_20_z_sink_wenable <= 0;
      _mul_20_z_sink_fifo_enq <= 0;
      __mul_20_stream_ivalid_1 <= 0;
      __mul_20_stream_ivalid_2 <= 0;
      __mul_20_stream_ivalid_3 <= 0;
      __mul_20_stream_ivalid_4 <= 0;
      __mul_20_stream_ivalid_5 <= 0;
      __mul_20_stream_ivalid_6 <= 0;
      __mul_20_stream_ivalid_7 <= 0;
      __mul_20_stream_ivalid_8 <= 0;
      _greaterthan_data_431 <= 0;
      _minus_data_433 <= 0;
      _greatereq_data_444 <= 0;
      __delay_data_1848__variable_428 <= 0;
      __delay_data_1851__variable_429 <= 0;
      __delay_data_1854__variable_430 <= 0;
      _sll_data_435 <= 0;
      __delay_data_1845_greaterthan_431 <= 0;
      __delay_data_1846_greatereq_444 <= 0;
      __delay_data_1849__delay_1848__variable_428 <= 0;
      __delay_data_1852__delay_1851__variable_429 <= 0;
      __delay_data_1855__delay_1854__variable_430 <= 0;
      _cond_data_441 <= 0;
      __delay_data_1847__delay_1846_greatereq_444 <= 0;
      __delay_data_1850__delay_1849__delay_1848__variable_428 <= 0;
      __delay_data_1853__delay_1852__delay_1851__variable_429 <= 0;
      __delay_data_1856__delay_1855__delay_1854__variable_430 <= 0;
      __muladd_madd_odata_reg_447 <= 0;
      __delay_data_1857__delay_1856__delay_1855____variable_430 <= 0;
      __delay_data_1858__delay_1857__delay_1856____variable_430 <= 0;
      __delay_data_1859__delay_1858__delay_1857____variable_430 <= 0;
      __delay_data_1860__delay_1859__delay_1858____variable_430 <= 0;
      _sra_data_448 <= 0;
      __variable_wdata_428 <= 0;
      __variable_wdata_429 <= 0;
      __variable_wdata_430 <= 0;
      _tmp_896 <= 0;
      _tmp_897 <= 0;
      _tmp_898 <= 0;
      _tmp_899 <= 0;
      _tmp_900 <= 0;
      _tmp_901 <= 0;
      _tmp_902 <= 0;
      _tmp_903 <= 0;
      _tmp_904 <= 0;
      _tmp_905 <= 0;
      _tmp_906 <= 0;
      _tmp_907 <= 0;
      _tmp_908 <= 0;
      _tmp_909 <= 0;
      _tmp_910 <= 0;
      _tmp_911 <= 0;
      _tmp_912 <= 0;
      _tmp_913 <= 0;
      _tmp_914 <= 0;
      _tmp_915 <= 0;
      _tmp_916 <= 0;
      _tmp_917 <= 0;
      _tmp_918 <= 0;
      _tmp_919 <= 0;
      _tmp_920 <= 0;
      _tmp_921 <= 0;
      _tmp_922 <= 0;
      _tmp_923 <= 0;
      _tmp_924 <= 0;
      _tmp_925 <= 0;
      _tmp_926 <= 0;
      _tmp_927 <= 0;
      _tmp_928 <= 0;
      _tmp_929 <= 0;
      _mul_20_busy_reg <= 0;
    end else begin
      if(_mul_20_stream_oready) begin
        _mul_20_x_source_ram_renable <= 0;
        _mul_20_x_source_fifo_deq <= 0;
      end 
      _mul_20_x_idle <= _mul_20_x_idle;
      if(_mul_20_stream_oready) begin
        _mul_20_y_source_ram_renable <= 0;
        _mul_20_y_source_fifo_deq <= 0;
      end 
      _mul_20_y_idle <= _mul_20_y_idle;
      if(_mul_20_stream_oready) begin
        _mul_20_rshift_source_ram_renable <= 0;
        _mul_20_rshift_source_fifo_deq <= 0;
      end 
      _mul_20_rshift_idle <= _mul_20_rshift_idle;
      if(_mul_20_stream_oready) begin
        _mul_20_z_sink_wenable <= 0;
        _mul_20_z_sink_fifo_enq <= 0;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_1 <= _mul_20_stream_ivalid;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_2 <= __mul_20_stream_ivalid_1;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_3 <= __mul_20_stream_ivalid_2;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_4 <= __mul_20_stream_ivalid_3;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_5 <= __mul_20_stream_ivalid_4;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_6 <= __mul_20_stream_ivalid_5;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_7 <= __mul_20_stream_ivalid_6;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_8 <= __mul_20_stream_ivalid_7;
      end 
      if(_mul_20_stream_oready) begin
        _greaterthan_data_431 <= mul_20_rshift_data > 1'sd0;
      end 
      if(_mul_20_stream_oready) begin
        _minus_data_433 <= mul_20_rshift_data - 2'sd1;
      end 
      if(_mul_20_stream_oready) begin
        _greatereq_data_444 <= mul_20_x_data >= 1'sd0;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1848__variable_428 <= mul_20_x_data;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1851__variable_429 <= mul_20_y_data;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1854__variable_430 <= mul_20_rshift_data;
      end 
      if(_mul_20_stream_oready) begin
        _sll_data_435 <= 2'sd1 << _minus_data_433;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1845_greaterthan_431 <= _greaterthan_data_431;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1846_greatereq_444 <= _greatereq_data_444;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1849__delay_1848__variable_428 <= __delay_data_1848__variable_428;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1852__delay_1851__variable_429 <= __delay_data_1851__variable_429;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1855__delay_1854__variable_430 <= __delay_data_1854__variable_430;
      end 
      if(_mul_20_stream_oready) begin
        _cond_data_441 <= (__delay_data_1845_greaterthan_431)? _sll_data_435 : 1'sd0;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1847__delay_1846_greatereq_444 <= __delay_data_1846_greatereq_444;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1850__delay_1849__delay_1848__variable_428 <= __delay_data_1849__delay_1848__variable_428;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1853__delay_1852__delay_1851__variable_429 <= __delay_data_1852__delay_1851__variable_429;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1856__delay_1855__delay_1854__variable_430 <= __delay_data_1855__delay_1854__variable_430;
      end 
      if(_mul_20_stream_oready) begin
        __muladd_madd_odata_reg_447 <= __muladd_madd_odata_447;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1857__delay_1856__delay_1855____variable_430 <= __delay_data_1856__delay_1855__delay_1854__variable_430;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1858__delay_1857__delay_1856____variable_430 <= __delay_data_1857__delay_1856__delay_1855____variable_430;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1859__delay_1858__delay_1857____variable_430 <= __delay_data_1858__delay_1857__delay_1856____variable_430;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1860__delay_1859__delay_1858____variable_430 <= __delay_data_1859__delay_1858__delay_1857____variable_430;
      end 
      if(_mul_20_stream_oready) begin
        _sra_data_448 <= __muladd_data_447 >>> __delay_data_1860__delay_1859__delay_1858____variable_430;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_428 <= _cond_data_1776;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_429 <= _cond_data_1443;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_430 <= __delay_data_2722__delay_2721_plus_1861;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_896 <= _mul_20_source_start;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_897 <= _tmp_896;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_898 <= _tmp_897;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_899 <= _mul_20_source_start;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_900 <= _tmp_899;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_901 <= _tmp_900;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_902 <= _tmp_901;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_903 <= _tmp_902;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_904 <= _tmp_903;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_905 <= _tmp_904;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_906 <= _tmp_905;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_907 <= _tmp_906;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_908 <= _tmp_907;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_909 <= _mul_20_source_stop;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_910 <= _tmp_909;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_911 <= _tmp_910;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_912 <= _tmp_911;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_913 <= _tmp_912;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_914 <= _tmp_913;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_915 <= _tmp_914;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_916 <= _tmp_915;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_917 <= _tmp_916;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_918 <= _tmp_917;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_919 <= _mul_20_source_busy;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_920 <= _tmp_919;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_921 <= _tmp_920;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_922 <= _tmp_921;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_923 <= _tmp_922;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_924 <= _tmp_923;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_925 <= _tmp_924;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_926 <= _tmp_925;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_927 <= _tmp_926;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_928 <= _tmp_927;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_929 <= _mul_20_sink_busy;
      end 
      if(!_mul_20_sink_busy && _tmp_929) begin
        _mul_20_busy_reg <= 0;
      end 
      if(_mul_20_source_busy) begin
        _mul_20_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_20_fsm_1 = 1;
  localparam _mul_20_fsm_2 = 2;
  localparam _mul_20_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_20_fsm <= _mul_20_fsm_init;
      _mul_20_source_start <= 0;
      _mul_20_source_busy <= 0;
      _mul_20_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_20_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_20_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_20_stream_oready && _tmp_898) begin
        _mul_20_stream_ivalid <= 1;
      end 
      if(_mul_20_stream_oready && 1'd0) begin
        _mul_20_stream_ivalid <= 0;
      end 
      case(_mul_20_fsm)
        _mul_20_fsm_init: begin
          if(_mul_20_run_flag) begin
            _mul_20_source_start <= 1;
          end 
          if(_mul_20_run_flag) begin
            _mul_20_fsm <= _mul_20_fsm_1;
          end 
        end
        _mul_20_fsm_1: begin
          if(_mul_20_source_start && _mul_20_stream_oready) begin
            _mul_20_source_start <= 0;
            _mul_20_source_busy <= 1;
          end 
          if(_mul_20_source_start && _mul_20_stream_oready) begin
            _mul_20_fsm <= _mul_20_fsm_2;
          end 
        end
        _mul_20_fsm_2: begin
          if(_mul_20_stream_oready) begin
            _mul_20_fsm <= _mul_20_fsm_3;
          end 
        end
        _mul_20_fsm_3: begin
          if(_mul_20_stream_oready && 1'd0) begin
            _mul_20_source_busy <= 0;
          end 
          if(_mul_20_stream_oready && 1'd0 && _mul_20_run_flag) begin
            _mul_20_source_start <= 1;
          end 
          if(_mul_20_stream_oready && 1'd0) begin
            _mul_20_fsm <= _mul_20_fsm_init;
          end 
          if(_mul_20_stream_oready && 1'd0 && _mul_20_run_flag) begin
            _mul_20_fsm <= _mul_20_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_21_x_source_ram_renable <= 0;
      _mul_21_x_source_fifo_deq <= 0;
      _mul_21_x_idle <= 1;
      _mul_21_y_source_ram_renable <= 0;
      _mul_21_y_source_fifo_deq <= 0;
      _mul_21_y_idle <= 1;
      _mul_21_rshift_source_ram_renable <= 0;
      _mul_21_rshift_source_fifo_deq <= 0;
      _mul_21_rshift_idle <= 1;
      _mul_21_z_sink_wenable <= 0;
      _mul_21_z_sink_fifo_enq <= 0;
      __mul_21_stream_ivalid_1 <= 0;
      __mul_21_stream_ivalid_2 <= 0;
      __mul_21_stream_ivalid_3 <= 0;
      __mul_21_stream_ivalid_4 <= 0;
      __mul_21_stream_ivalid_5 <= 0;
      __mul_21_stream_ivalid_6 <= 0;
      __mul_21_stream_ivalid_7 <= 0;
      __mul_21_stream_ivalid_8 <= 0;
      _greaterthan_data_452 <= 0;
      _minus_data_454 <= 0;
      _greatereq_data_465 <= 0;
      __delay_data_1867__variable_449 <= 0;
      __delay_data_1870__variable_450 <= 0;
      __delay_data_1873__variable_451 <= 0;
      _sll_data_456 <= 0;
      __delay_data_1864_greaterthan_452 <= 0;
      __delay_data_1865_greatereq_465 <= 0;
      __delay_data_1868__delay_1867__variable_449 <= 0;
      __delay_data_1871__delay_1870__variable_450 <= 0;
      __delay_data_1874__delay_1873__variable_451 <= 0;
      _cond_data_462 <= 0;
      __delay_data_1866__delay_1865_greatereq_465 <= 0;
      __delay_data_1869__delay_1868__delay_1867__variable_449 <= 0;
      __delay_data_1872__delay_1871__delay_1870__variable_450 <= 0;
      __delay_data_1875__delay_1874__delay_1873__variable_451 <= 0;
      __muladd_madd_odata_reg_468 <= 0;
      __delay_data_1876__delay_1875__delay_1874____variable_451 <= 0;
      __delay_data_1877__delay_1876__delay_1875____variable_451 <= 0;
      __delay_data_1878__delay_1877__delay_1876____variable_451 <= 0;
      __delay_data_1879__delay_1878__delay_1877____variable_451 <= 0;
      _sra_data_469 <= 0;
      __variable_wdata_449 <= 0;
      __variable_wdata_450 <= 0;
      __variable_wdata_451 <= 0;
      _tmp_930 <= 0;
      _tmp_931 <= 0;
      _tmp_932 <= 0;
      _tmp_933 <= 0;
      _tmp_934 <= 0;
      _tmp_935 <= 0;
      _tmp_936 <= 0;
      _tmp_937 <= 0;
      _tmp_938 <= 0;
      _tmp_939 <= 0;
      _tmp_940 <= 0;
      _tmp_941 <= 0;
      _tmp_942 <= 0;
      _tmp_943 <= 0;
      _tmp_944 <= 0;
      _tmp_945 <= 0;
      _tmp_946 <= 0;
      _tmp_947 <= 0;
      _tmp_948 <= 0;
      _tmp_949 <= 0;
      _tmp_950 <= 0;
      _tmp_951 <= 0;
      _tmp_952 <= 0;
      _tmp_953 <= 0;
      _tmp_954 <= 0;
      _tmp_955 <= 0;
      _tmp_956 <= 0;
      _tmp_957 <= 0;
      _tmp_958 <= 0;
      _tmp_959 <= 0;
      _tmp_960 <= 0;
      _tmp_961 <= 0;
      _tmp_962 <= 0;
      _tmp_963 <= 0;
      _mul_21_busy_reg <= 0;
    end else begin
      if(_mul_21_stream_oready) begin
        _mul_21_x_source_ram_renable <= 0;
        _mul_21_x_source_fifo_deq <= 0;
      end 
      _mul_21_x_idle <= _mul_21_x_idle;
      if(_mul_21_stream_oready) begin
        _mul_21_y_source_ram_renable <= 0;
        _mul_21_y_source_fifo_deq <= 0;
      end 
      _mul_21_y_idle <= _mul_21_y_idle;
      if(_mul_21_stream_oready) begin
        _mul_21_rshift_source_ram_renable <= 0;
        _mul_21_rshift_source_fifo_deq <= 0;
      end 
      _mul_21_rshift_idle <= _mul_21_rshift_idle;
      if(_mul_21_stream_oready) begin
        _mul_21_z_sink_wenable <= 0;
        _mul_21_z_sink_fifo_enq <= 0;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_1 <= _mul_21_stream_ivalid;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_2 <= __mul_21_stream_ivalid_1;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_3 <= __mul_21_stream_ivalid_2;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_4 <= __mul_21_stream_ivalid_3;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_5 <= __mul_21_stream_ivalid_4;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_6 <= __mul_21_stream_ivalid_5;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_7 <= __mul_21_stream_ivalid_6;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_8 <= __mul_21_stream_ivalid_7;
      end 
      if(_mul_21_stream_oready) begin
        _greaterthan_data_452 <= mul_21_rshift_data > 1'sd0;
      end 
      if(_mul_21_stream_oready) begin
        _minus_data_454 <= mul_21_rshift_data - 2'sd1;
      end 
      if(_mul_21_stream_oready) begin
        _greatereq_data_465 <= mul_21_x_data >= 1'sd0;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1867__variable_449 <= mul_21_x_data;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1870__variable_450 <= mul_21_y_data;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1873__variable_451 <= mul_21_rshift_data;
      end 
      if(_mul_21_stream_oready) begin
        _sll_data_456 <= 2'sd1 << _minus_data_454;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1864_greaterthan_452 <= _greaterthan_data_452;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1865_greatereq_465 <= _greatereq_data_465;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1868__delay_1867__variable_449 <= __delay_data_1867__variable_449;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1871__delay_1870__variable_450 <= __delay_data_1870__variable_450;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1874__delay_1873__variable_451 <= __delay_data_1873__variable_451;
      end 
      if(_mul_21_stream_oready) begin
        _cond_data_462 <= (__delay_data_1864_greaterthan_452)? _sll_data_456 : 1'sd0;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1866__delay_1865_greatereq_465 <= __delay_data_1865_greatereq_465;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1869__delay_1868__delay_1867__variable_449 <= __delay_data_1868__delay_1867__variable_449;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1872__delay_1871__delay_1870__variable_450 <= __delay_data_1871__delay_1870__variable_450;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1875__delay_1874__delay_1873__variable_451 <= __delay_data_1874__delay_1873__variable_451;
      end 
      if(_mul_21_stream_oready) begin
        __muladd_madd_odata_reg_468 <= __muladd_madd_odata_468;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1876__delay_1875__delay_1874____variable_451 <= __delay_data_1875__delay_1874__delay_1873__variable_451;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1877__delay_1876__delay_1875____variable_451 <= __delay_data_1876__delay_1875__delay_1874____variable_451;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1878__delay_1877__delay_1876____variable_451 <= __delay_data_1877__delay_1876__delay_1875____variable_451;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1879__delay_1878__delay_1877____variable_451 <= __delay_data_1878__delay_1877__delay_1876____variable_451;
      end 
      if(_mul_21_stream_oready) begin
        _sra_data_469 <= __muladd_data_468 >>> __delay_data_1879__delay_1878__delay_1877____variable_451;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_449 <= _cond_data_1778;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_450 <= _cond_data_1445;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_451 <= __delay_data_2739__delay_2738_plus_1880;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_930 <= _mul_21_source_start;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_931 <= _tmp_930;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_932 <= _tmp_931;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_933 <= _mul_21_source_start;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_934 <= _tmp_933;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_935 <= _tmp_934;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_936 <= _tmp_935;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_937 <= _tmp_936;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_938 <= _tmp_937;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_939 <= _tmp_938;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_940 <= _tmp_939;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_941 <= _tmp_940;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_942 <= _tmp_941;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_943 <= _mul_21_source_stop;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_944 <= _tmp_943;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_945 <= _tmp_944;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_946 <= _tmp_945;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_947 <= _tmp_946;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_948 <= _tmp_947;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_949 <= _tmp_948;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_950 <= _tmp_949;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_951 <= _tmp_950;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_952 <= _tmp_951;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_953 <= _mul_21_source_busy;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_954 <= _tmp_953;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_955 <= _tmp_954;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_956 <= _tmp_955;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_957 <= _tmp_956;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_958 <= _tmp_957;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_959 <= _tmp_958;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_960 <= _tmp_959;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_961 <= _tmp_960;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_962 <= _tmp_961;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_963 <= _mul_21_sink_busy;
      end 
      if(!_mul_21_sink_busy && _tmp_963) begin
        _mul_21_busy_reg <= 0;
      end 
      if(_mul_21_source_busy) begin
        _mul_21_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_21_fsm_1 = 1;
  localparam _mul_21_fsm_2 = 2;
  localparam _mul_21_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_21_fsm <= _mul_21_fsm_init;
      _mul_21_source_start <= 0;
      _mul_21_source_busy <= 0;
      _mul_21_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_21_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_21_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_21_stream_oready && _tmp_932) begin
        _mul_21_stream_ivalid <= 1;
      end 
      if(_mul_21_stream_oready && 1'd0) begin
        _mul_21_stream_ivalid <= 0;
      end 
      case(_mul_21_fsm)
        _mul_21_fsm_init: begin
          if(_mul_21_run_flag) begin
            _mul_21_source_start <= 1;
          end 
          if(_mul_21_run_flag) begin
            _mul_21_fsm <= _mul_21_fsm_1;
          end 
        end
        _mul_21_fsm_1: begin
          if(_mul_21_source_start && _mul_21_stream_oready) begin
            _mul_21_source_start <= 0;
            _mul_21_source_busy <= 1;
          end 
          if(_mul_21_source_start && _mul_21_stream_oready) begin
            _mul_21_fsm <= _mul_21_fsm_2;
          end 
        end
        _mul_21_fsm_2: begin
          if(_mul_21_stream_oready) begin
            _mul_21_fsm <= _mul_21_fsm_3;
          end 
        end
        _mul_21_fsm_3: begin
          if(_mul_21_stream_oready && 1'd0) begin
            _mul_21_source_busy <= 0;
          end 
          if(_mul_21_stream_oready && 1'd0 && _mul_21_run_flag) begin
            _mul_21_source_start <= 1;
          end 
          if(_mul_21_stream_oready && 1'd0) begin
            _mul_21_fsm <= _mul_21_fsm_init;
          end 
          if(_mul_21_stream_oready && 1'd0 && _mul_21_run_flag) begin
            _mul_21_fsm <= _mul_21_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_22_x_source_ram_renable <= 0;
      _mul_22_x_source_fifo_deq <= 0;
      _mul_22_x_idle <= 1;
      _mul_22_y_source_ram_renable <= 0;
      _mul_22_y_source_fifo_deq <= 0;
      _mul_22_y_idle <= 1;
      _mul_22_rshift_source_ram_renable <= 0;
      _mul_22_rshift_source_fifo_deq <= 0;
      _mul_22_rshift_idle <= 1;
      _mul_22_z_sink_wenable <= 0;
      _mul_22_z_sink_fifo_enq <= 0;
      __mul_22_stream_ivalid_1 <= 0;
      __mul_22_stream_ivalid_2 <= 0;
      __mul_22_stream_ivalid_3 <= 0;
      __mul_22_stream_ivalid_4 <= 0;
      __mul_22_stream_ivalid_5 <= 0;
      __mul_22_stream_ivalid_6 <= 0;
      __mul_22_stream_ivalid_7 <= 0;
      __mul_22_stream_ivalid_8 <= 0;
      _greaterthan_data_473 <= 0;
      _minus_data_475 <= 0;
      _greatereq_data_486 <= 0;
      __delay_data_1886__variable_470 <= 0;
      __delay_data_1889__variable_471 <= 0;
      __delay_data_1892__variable_472 <= 0;
      _sll_data_477 <= 0;
      __delay_data_1883_greaterthan_473 <= 0;
      __delay_data_1884_greatereq_486 <= 0;
      __delay_data_1887__delay_1886__variable_470 <= 0;
      __delay_data_1890__delay_1889__variable_471 <= 0;
      __delay_data_1893__delay_1892__variable_472 <= 0;
      _cond_data_483 <= 0;
      __delay_data_1885__delay_1884_greatereq_486 <= 0;
      __delay_data_1888__delay_1887__delay_1886__variable_470 <= 0;
      __delay_data_1891__delay_1890__delay_1889__variable_471 <= 0;
      __delay_data_1894__delay_1893__delay_1892__variable_472 <= 0;
      __muladd_madd_odata_reg_489 <= 0;
      __delay_data_1895__delay_1894__delay_1893____variable_472 <= 0;
      __delay_data_1896__delay_1895__delay_1894____variable_472 <= 0;
      __delay_data_1897__delay_1896__delay_1895____variable_472 <= 0;
      __delay_data_1898__delay_1897__delay_1896____variable_472 <= 0;
      _sra_data_490 <= 0;
      __variable_wdata_470 <= 0;
      __variable_wdata_471 <= 0;
      __variable_wdata_472 <= 0;
      _tmp_964 <= 0;
      _tmp_965 <= 0;
      _tmp_966 <= 0;
      _tmp_967 <= 0;
      _tmp_968 <= 0;
      _tmp_969 <= 0;
      _tmp_970 <= 0;
      _tmp_971 <= 0;
      _tmp_972 <= 0;
      _tmp_973 <= 0;
      _tmp_974 <= 0;
      _tmp_975 <= 0;
      _tmp_976 <= 0;
      _tmp_977 <= 0;
      _tmp_978 <= 0;
      _tmp_979 <= 0;
      _tmp_980 <= 0;
      _tmp_981 <= 0;
      _tmp_982 <= 0;
      _tmp_983 <= 0;
      _tmp_984 <= 0;
      _tmp_985 <= 0;
      _tmp_986 <= 0;
      _tmp_987 <= 0;
      _tmp_988 <= 0;
      _tmp_989 <= 0;
      _tmp_990 <= 0;
      _tmp_991 <= 0;
      _tmp_992 <= 0;
      _tmp_993 <= 0;
      _tmp_994 <= 0;
      _tmp_995 <= 0;
      _tmp_996 <= 0;
      _tmp_997 <= 0;
      _mul_22_busy_reg <= 0;
    end else begin
      if(_mul_22_stream_oready) begin
        _mul_22_x_source_ram_renable <= 0;
        _mul_22_x_source_fifo_deq <= 0;
      end 
      _mul_22_x_idle <= _mul_22_x_idle;
      if(_mul_22_stream_oready) begin
        _mul_22_y_source_ram_renable <= 0;
        _mul_22_y_source_fifo_deq <= 0;
      end 
      _mul_22_y_idle <= _mul_22_y_idle;
      if(_mul_22_stream_oready) begin
        _mul_22_rshift_source_ram_renable <= 0;
        _mul_22_rshift_source_fifo_deq <= 0;
      end 
      _mul_22_rshift_idle <= _mul_22_rshift_idle;
      if(_mul_22_stream_oready) begin
        _mul_22_z_sink_wenable <= 0;
        _mul_22_z_sink_fifo_enq <= 0;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_1 <= _mul_22_stream_ivalid;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_2 <= __mul_22_stream_ivalid_1;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_3 <= __mul_22_stream_ivalid_2;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_4 <= __mul_22_stream_ivalid_3;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_5 <= __mul_22_stream_ivalid_4;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_6 <= __mul_22_stream_ivalid_5;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_7 <= __mul_22_stream_ivalid_6;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_8 <= __mul_22_stream_ivalid_7;
      end 
      if(_mul_22_stream_oready) begin
        _greaterthan_data_473 <= mul_22_rshift_data > 1'sd0;
      end 
      if(_mul_22_stream_oready) begin
        _minus_data_475 <= mul_22_rshift_data - 2'sd1;
      end 
      if(_mul_22_stream_oready) begin
        _greatereq_data_486 <= mul_22_x_data >= 1'sd0;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1886__variable_470 <= mul_22_x_data;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1889__variable_471 <= mul_22_y_data;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1892__variable_472 <= mul_22_rshift_data;
      end 
      if(_mul_22_stream_oready) begin
        _sll_data_477 <= 2'sd1 << _minus_data_475;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1883_greaterthan_473 <= _greaterthan_data_473;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1884_greatereq_486 <= _greatereq_data_486;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1887__delay_1886__variable_470 <= __delay_data_1886__variable_470;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1890__delay_1889__variable_471 <= __delay_data_1889__variable_471;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1893__delay_1892__variable_472 <= __delay_data_1892__variable_472;
      end 
      if(_mul_22_stream_oready) begin
        _cond_data_483 <= (__delay_data_1883_greaterthan_473)? _sll_data_477 : 1'sd0;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1885__delay_1884_greatereq_486 <= __delay_data_1884_greatereq_486;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1888__delay_1887__delay_1886__variable_470 <= __delay_data_1887__delay_1886__variable_470;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1891__delay_1890__delay_1889__variable_471 <= __delay_data_1890__delay_1889__variable_471;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1894__delay_1893__delay_1892__variable_472 <= __delay_data_1893__delay_1892__variable_472;
      end 
      if(_mul_22_stream_oready) begin
        __muladd_madd_odata_reg_489 <= __muladd_madd_odata_489;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1895__delay_1894__delay_1893____variable_472 <= __delay_data_1894__delay_1893__delay_1892__variable_472;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1896__delay_1895__delay_1894____variable_472 <= __delay_data_1895__delay_1894__delay_1893____variable_472;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1897__delay_1896__delay_1895____variable_472 <= __delay_data_1896__delay_1895__delay_1894____variable_472;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_1898__delay_1897__delay_1896____variable_472 <= __delay_data_1897__delay_1896__delay_1895____variable_472;
      end 
      if(_mul_22_stream_oready) begin
        _sra_data_490 <= __muladd_data_489 >>> __delay_data_1898__delay_1897__delay_1896____variable_472;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_470 <= _cond_data_1780;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_471 <= _cond_data_1447;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_472 <= __delay_data_2756__delay_2755_plus_1899;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_964 <= _mul_22_source_start;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_965 <= _tmp_964;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_966 <= _tmp_965;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_967 <= _mul_22_source_start;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_968 <= _tmp_967;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_969 <= _tmp_968;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_970 <= _tmp_969;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_971 <= _tmp_970;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_972 <= _tmp_971;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_973 <= _tmp_972;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_974 <= _tmp_973;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_975 <= _tmp_974;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_976 <= _tmp_975;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_977 <= _mul_22_source_stop;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_978 <= _tmp_977;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_979 <= _tmp_978;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_980 <= _tmp_979;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_981 <= _tmp_980;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_982 <= _tmp_981;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_983 <= _tmp_982;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_984 <= _tmp_983;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_985 <= _tmp_984;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_986 <= _tmp_985;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_987 <= _mul_22_source_busy;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_988 <= _tmp_987;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_989 <= _tmp_988;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_990 <= _tmp_989;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_991 <= _tmp_990;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_992 <= _tmp_991;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_993 <= _tmp_992;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_994 <= _tmp_993;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_995 <= _tmp_994;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_996 <= _tmp_995;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_997 <= _mul_22_sink_busy;
      end 
      if(!_mul_22_sink_busy && _tmp_997) begin
        _mul_22_busy_reg <= 0;
      end 
      if(_mul_22_source_busy) begin
        _mul_22_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_22_fsm_1 = 1;
  localparam _mul_22_fsm_2 = 2;
  localparam _mul_22_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_22_fsm <= _mul_22_fsm_init;
      _mul_22_source_start <= 0;
      _mul_22_source_busy <= 0;
      _mul_22_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_22_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_22_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_22_stream_oready && _tmp_966) begin
        _mul_22_stream_ivalid <= 1;
      end 
      if(_mul_22_stream_oready && 1'd0) begin
        _mul_22_stream_ivalid <= 0;
      end 
      case(_mul_22_fsm)
        _mul_22_fsm_init: begin
          if(_mul_22_run_flag) begin
            _mul_22_source_start <= 1;
          end 
          if(_mul_22_run_flag) begin
            _mul_22_fsm <= _mul_22_fsm_1;
          end 
        end
        _mul_22_fsm_1: begin
          if(_mul_22_source_start && _mul_22_stream_oready) begin
            _mul_22_source_start <= 0;
            _mul_22_source_busy <= 1;
          end 
          if(_mul_22_source_start && _mul_22_stream_oready) begin
            _mul_22_fsm <= _mul_22_fsm_2;
          end 
        end
        _mul_22_fsm_2: begin
          if(_mul_22_stream_oready) begin
            _mul_22_fsm <= _mul_22_fsm_3;
          end 
        end
        _mul_22_fsm_3: begin
          if(_mul_22_stream_oready && 1'd0) begin
            _mul_22_source_busy <= 0;
          end 
          if(_mul_22_stream_oready && 1'd0 && _mul_22_run_flag) begin
            _mul_22_source_start <= 1;
          end 
          if(_mul_22_stream_oready && 1'd0) begin
            _mul_22_fsm <= _mul_22_fsm_init;
          end 
          if(_mul_22_stream_oready && 1'd0 && _mul_22_run_flag) begin
            _mul_22_fsm <= _mul_22_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_23_x_source_ram_renable <= 0;
      _mul_23_x_source_fifo_deq <= 0;
      _mul_23_x_idle <= 1;
      _mul_23_y_source_ram_renable <= 0;
      _mul_23_y_source_fifo_deq <= 0;
      _mul_23_y_idle <= 1;
      _mul_23_rshift_source_ram_renable <= 0;
      _mul_23_rshift_source_fifo_deq <= 0;
      _mul_23_rshift_idle <= 1;
      _mul_23_z_sink_wenable <= 0;
      _mul_23_z_sink_fifo_enq <= 0;
      __mul_23_stream_ivalid_1 <= 0;
      __mul_23_stream_ivalid_2 <= 0;
      __mul_23_stream_ivalid_3 <= 0;
      __mul_23_stream_ivalid_4 <= 0;
      __mul_23_stream_ivalid_5 <= 0;
      __mul_23_stream_ivalid_6 <= 0;
      __mul_23_stream_ivalid_7 <= 0;
      __mul_23_stream_ivalid_8 <= 0;
      _greaterthan_data_494 <= 0;
      _minus_data_496 <= 0;
      _greatereq_data_507 <= 0;
      __delay_data_1905__variable_491 <= 0;
      __delay_data_1908__variable_492 <= 0;
      __delay_data_1911__variable_493 <= 0;
      _sll_data_498 <= 0;
      __delay_data_1902_greaterthan_494 <= 0;
      __delay_data_1903_greatereq_507 <= 0;
      __delay_data_1906__delay_1905__variable_491 <= 0;
      __delay_data_1909__delay_1908__variable_492 <= 0;
      __delay_data_1912__delay_1911__variable_493 <= 0;
      _cond_data_504 <= 0;
      __delay_data_1904__delay_1903_greatereq_507 <= 0;
      __delay_data_1907__delay_1906__delay_1905__variable_491 <= 0;
      __delay_data_1910__delay_1909__delay_1908__variable_492 <= 0;
      __delay_data_1913__delay_1912__delay_1911__variable_493 <= 0;
      __muladd_madd_odata_reg_510 <= 0;
      __delay_data_1914__delay_1913__delay_1912____variable_493 <= 0;
      __delay_data_1915__delay_1914__delay_1913____variable_493 <= 0;
      __delay_data_1916__delay_1915__delay_1914____variable_493 <= 0;
      __delay_data_1917__delay_1916__delay_1915____variable_493 <= 0;
      _sra_data_511 <= 0;
      __variable_wdata_491 <= 0;
      __variable_wdata_492 <= 0;
      __variable_wdata_493 <= 0;
      _tmp_998 <= 0;
      _tmp_999 <= 0;
      _tmp_1000 <= 0;
      _tmp_1001 <= 0;
      _tmp_1002 <= 0;
      _tmp_1003 <= 0;
      _tmp_1004 <= 0;
      _tmp_1005 <= 0;
      _tmp_1006 <= 0;
      _tmp_1007 <= 0;
      _tmp_1008 <= 0;
      _tmp_1009 <= 0;
      _tmp_1010 <= 0;
      _tmp_1011 <= 0;
      _tmp_1012 <= 0;
      _tmp_1013 <= 0;
      _tmp_1014 <= 0;
      _tmp_1015 <= 0;
      _tmp_1016 <= 0;
      _tmp_1017 <= 0;
      _tmp_1018 <= 0;
      _tmp_1019 <= 0;
      _tmp_1020 <= 0;
      _tmp_1021 <= 0;
      _tmp_1022 <= 0;
      _tmp_1023 <= 0;
      _tmp_1024 <= 0;
      _tmp_1025 <= 0;
      _tmp_1026 <= 0;
      _tmp_1027 <= 0;
      _tmp_1028 <= 0;
      _tmp_1029 <= 0;
      _tmp_1030 <= 0;
      _tmp_1031 <= 0;
      _mul_23_busy_reg <= 0;
    end else begin
      if(_mul_23_stream_oready) begin
        _mul_23_x_source_ram_renable <= 0;
        _mul_23_x_source_fifo_deq <= 0;
      end 
      _mul_23_x_idle <= _mul_23_x_idle;
      if(_mul_23_stream_oready) begin
        _mul_23_y_source_ram_renable <= 0;
        _mul_23_y_source_fifo_deq <= 0;
      end 
      _mul_23_y_idle <= _mul_23_y_idle;
      if(_mul_23_stream_oready) begin
        _mul_23_rshift_source_ram_renable <= 0;
        _mul_23_rshift_source_fifo_deq <= 0;
      end 
      _mul_23_rshift_idle <= _mul_23_rshift_idle;
      if(_mul_23_stream_oready) begin
        _mul_23_z_sink_wenable <= 0;
        _mul_23_z_sink_fifo_enq <= 0;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_1 <= _mul_23_stream_ivalid;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_2 <= __mul_23_stream_ivalid_1;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_3 <= __mul_23_stream_ivalid_2;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_4 <= __mul_23_stream_ivalid_3;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_5 <= __mul_23_stream_ivalid_4;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_6 <= __mul_23_stream_ivalid_5;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_7 <= __mul_23_stream_ivalid_6;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_8 <= __mul_23_stream_ivalid_7;
      end 
      if(_mul_23_stream_oready) begin
        _greaterthan_data_494 <= mul_23_rshift_data > 1'sd0;
      end 
      if(_mul_23_stream_oready) begin
        _minus_data_496 <= mul_23_rshift_data - 2'sd1;
      end 
      if(_mul_23_stream_oready) begin
        _greatereq_data_507 <= mul_23_x_data >= 1'sd0;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1905__variable_491 <= mul_23_x_data;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1908__variable_492 <= mul_23_y_data;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1911__variable_493 <= mul_23_rshift_data;
      end 
      if(_mul_23_stream_oready) begin
        _sll_data_498 <= 2'sd1 << _minus_data_496;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1902_greaterthan_494 <= _greaterthan_data_494;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1903_greatereq_507 <= _greatereq_data_507;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1906__delay_1905__variable_491 <= __delay_data_1905__variable_491;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1909__delay_1908__variable_492 <= __delay_data_1908__variable_492;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1912__delay_1911__variable_493 <= __delay_data_1911__variable_493;
      end 
      if(_mul_23_stream_oready) begin
        _cond_data_504 <= (__delay_data_1902_greaterthan_494)? _sll_data_498 : 1'sd0;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1904__delay_1903_greatereq_507 <= __delay_data_1903_greatereq_507;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1907__delay_1906__delay_1905__variable_491 <= __delay_data_1906__delay_1905__variable_491;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1910__delay_1909__delay_1908__variable_492 <= __delay_data_1909__delay_1908__variable_492;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1913__delay_1912__delay_1911__variable_493 <= __delay_data_1912__delay_1911__variable_493;
      end 
      if(_mul_23_stream_oready) begin
        __muladd_madd_odata_reg_510 <= __muladd_madd_odata_510;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1914__delay_1913__delay_1912____variable_493 <= __delay_data_1913__delay_1912__delay_1911__variable_493;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1915__delay_1914__delay_1913____variable_493 <= __delay_data_1914__delay_1913__delay_1912____variable_493;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1916__delay_1915__delay_1914____variable_493 <= __delay_data_1915__delay_1914__delay_1913____variable_493;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_1917__delay_1916__delay_1915____variable_493 <= __delay_data_1916__delay_1915__delay_1914____variable_493;
      end 
      if(_mul_23_stream_oready) begin
        _sra_data_511 <= __muladd_data_510 >>> __delay_data_1917__delay_1916__delay_1915____variable_493;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_491 <= _cond_data_1782;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_492 <= _cond_data_1449;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_493 <= __delay_data_2773__delay_2772_plus_1918;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_998 <= _mul_23_source_start;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_999 <= _tmp_998;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1000 <= _tmp_999;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1001 <= _mul_23_source_start;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1002 <= _tmp_1001;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1003 <= _tmp_1002;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1004 <= _tmp_1003;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1005 <= _tmp_1004;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1006 <= _tmp_1005;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1007 <= _tmp_1006;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1008 <= _tmp_1007;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1009 <= _tmp_1008;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1010 <= _tmp_1009;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1011 <= _mul_23_source_stop;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1012 <= _tmp_1011;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1013 <= _tmp_1012;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1014 <= _tmp_1013;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1015 <= _tmp_1014;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1016 <= _tmp_1015;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1017 <= _tmp_1016;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1018 <= _tmp_1017;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1019 <= _tmp_1018;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1020 <= _tmp_1019;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1021 <= _mul_23_source_busy;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1022 <= _tmp_1021;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1023 <= _tmp_1022;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1024 <= _tmp_1023;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1025 <= _tmp_1024;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1026 <= _tmp_1025;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1027 <= _tmp_1026;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1028 <= _tmp_1027;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1029 <= _tmp_1028;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1030 <= _tmp_1029;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_1031 <= _mul_23_sink_busy;
      end 
      if(!_mul_23_sink_busy && _tmp_1031) begin
        _mul_23_busy_reg <= 0;
      end 
      if(_mul_23_source_busy) begin
        _mul_23_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_23_fsm_1 = 1;
  localparam _mul_23_fsm_2 = 2;
  localparam _mul_23_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_23_fsm <= _mul_23_fsm_init;
      _mul_23_source_start <= 0;
      _mul_23_source_busy <= 0;
      _mul_23_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_23_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_23_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_23_stream_oready && _tmp_1000) begin
        _mul_23_stream_ivalid <= 1;
      end 
      if(_mul_23_stream_oready && 1'd0) begin
        _mul_23_stream_ivalid <= 0;
      end 
      case(_mul_23_fsm)
        _mul_23_fsm_init: begin
          if(_mul_23_run_flag) begin
            _mul_23_source_start <= 1;
          end 
          if(_mul_23_run_flag) begin
            _mul_23_fsm <= _mul_23_fsm_1;
          end 
        end
        _mul_23_fsm_1: begin
          if(_mul_23_source_start && _mul_23_stream_oready) begin
            _mul_23_source_start <= 0;
            _mul_23_source_busy <= 1;
          end 
          if(_mul_23_source_start && _mul_23_stream_oready) begin
            _mul_23_fsm <= _mul_23_fsm_2;
          end 
        end
        _mul_23_fsm_2: begin
          if(_mul_23_stream_oready) begin
            _mul_23_fsm <= _mul_23_fsm_3;
          end 
        end
        _mul_23_fsm_3: begin
          if(_mul_23_stream_oready && 1'd0) begin
            _mul_23_source_busy <= 0;
          end 
          if(_mul_23_stream_oready && 1'd0 && _mul_23_run_flag) begin
            _mul_23_source_start <= 1;
          end 
          if(_mul_23_stream_oready && 1'd0) begin
            _mul_23_fsm <= _mul_23_fsm_init;
          end 
          if(_mul_23_stream_oready && 1'd0 && _mul_23_run_flag) begin
            _mul_23_fsm <= _mul_23_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_24_x_source_ram_renable <= 0;
      _mul_24_x_source_fifo_deq <= 0;
      _mul_24_x_idle <= 1;
      _mul_24_y_source_ram_renable <= 0;
      _mul_24_y_source_fifo_deq <= 0;
      _mul_24_y_idle <= 1;
      _mul_24_rshift_source_ram_renable <= 0;
      _mul_24_rshift_source_fifo_deq <= 0;
      _mul_24_rshift_idle <= 1;
      _mul_24_z_sink_wenable <= 0;
      _mul_24_z_sink_fifo_enq <= 0;
      __mul_24_stream_ivalid_1 <= 0;
      __mul_24_stream_ivalid_2 <= 0;
      __mul_24_stream_ivalid_3 <= 0;
      __mul_24_stream_ivalid_4 <= 0;
      __mul_24_stream_ivalid_5 <= 0;
      __mul_24_stream_ivalid_6 <= 0;
      __mul_24_stream_ivalid_7 <= 0;
      __mul_24_stream_ivalid_8 <= 0;
      _greaterthan_data_515 <= 0;
      _minus_data_517 <= 0;
      _greatereq_data_528 <= 0;
      __delay_data_1924__variable_512 <= 0;
      __delay_data_1927__variable_513 <= 0;
      __delay_data_1930__variable_514 <= 0;
      _sll_data_519 <= 0;
      __delay_data_1921_greaterthan_515 <= 0;
      __delay_data_1922_greatereq_528 <= 0;
      __delay_data_1925__delay_1924__variable_512 <= 0;
      __delay_data_1928__delay_1927__variable_513 <= 0;
      __delay_data_1931__delay_1930__variable_514 <= 0;
      _cond_data_525 <= 0;
      __delay_data_1923__delay_1922_greatereq_528 <= 0;
      __delay_data_1926__delay_1925__delay_1924__variable_512 <= 0;
      __delay_data_1929__delay_1928__delay_1927__variable_513 <= 0;
      __delay_data_1932__delay_1931__delay_1930__variable_514 <= 0;
      __muladd_madd_odata_reg_531 <= 0;
      __delay_data_1933__delay_1932__delay_1931____variable_514 <= 0;
      __delay_data_1934__delay_1933__delay_1932____variable_514 <= 0;
      __delay_data_1935__delay_1934__delay_1933____variable_514 <= 0;
      __delay_data_1936__delay_1935__delay_1934____variable_514 <= 0;
      _sra_data_532 <= 0;
      __variable_wdata_512 <= 0;
      __variable_wdata_513 <= 0;
      __variable_wdata_514 <= 0;
      _tmp_1032 <= 0;
      _tmp_1033 <= 0;
      _tmp_1034 <= 0;
      _tmp_1035 <= 0;
      _tmp_1036 <= 0;
      _tmp_1037 <= 0;
      _tmp_1038 <= 0;
      _tmp_1039 <= 0;
      _tmp_1040 <= 0;
      _tmp_1041 <= 0;
      _tmp_1042 <= 0;
      _tmp_1043 <= 0;
      _tmp_1044 <= 0;
      _tmp_1045 <= 0;
      _tmp_1046 <= 0;
      _tmp_1047 <= 0;
      _tmp_1048 <= 0;
      _tmp_1049 <= 0;
      _tmp_1050 <= 0;
      _tmp_1051 <= 0;
      _tmp_1052 <= 0;
      _tmp_1053 <= 0;
      _tmp_1054 <= 0;
      _tmp_1055 <= 0;
      _tmp_1056 <= 0;
      _tmp_1057 <= 0;
      _tmp_1058 <= 0;
      _tmp_1059 <= 0;
      _tmp_1060 <= 0;
      _tmp_1061 <= 0;
      _tmp_1062 <= 0;
      _tmp_1063 <= 0;
      _tmp_1064 <= 0;
      _tmp_1065 <= 0;
      _mul_24_busy_reg <= 0;
    end else begin
      if(_mul_24_stream_oready) begin
        _mul_24_x_source_ram_renable <= 0;
        _mul_24_x_source_fifo_deq <= 0;
      end 
      _mul_24_x_idle <= _mul_24_x_idle;
      if(_mul_24_stream_oready) begin
        _mul_24_y_source_ram_renable <= 0;
        _mul_24_y_source_fifo_deq <= 0;
      end 
      _mul_24_y_idle <= _mul_24_y_idle;
      if(_mul_24_stream_oready) begin
        _mul_24_rshift_source_ram_renable <= 0;
        _mul_24_rshift_source_fifo_deq <= 0;
      end 
      _mul_24_rshift_idle <= _mul_24_rshift_idle;
      if(_mul_24_stream_oready) begin
        _mul_24_z_sink_wenable <= 0;
        _mul_24_z_sink_fifo_enq <= 0;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_1 <= _mul_24_stream_ivalid;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_2 <= __mul_24_stream_ivalid_1;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_3 <= __mul_24_stream_ivalid_2;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_4 <= __mul_24_stream_ivalid_3;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_5 <= __mul_24_stream_ivalid_4;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_6 <= __mul_24_stream_ivalid_5;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_7 <= __mul_24_stream_ivalid_6;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_8 <= __mul_24_stream_ivalid_7;
      end 
      if(_mul_24_stream_oready) begin
        _greaterthan_data_515 <= mul_24_rshift_data > 1'sd0;
      end 
      if(_mul_24_stream_oready) begin
        _minus_data_517 <= mul_24_rshift_data - 2'sd1;
      end 
      if(_mul_24_stream_oready) begin
        _greatereq_data_528 <= mul_24_x_data >= 1'sd0;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1924__variable_512 <= mul_24_x_data;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1927__variable_513 <= mul_24_y_data;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1930__variable_514 <= mul_24_rshift_data;
      end 
      if(_mul_24_stream_oready) begin
        _sll_data_519 <= 2'sd1 << _minus_data_517;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1921_greaterthan_515 <= _greaterthan_data_515;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1922_greatereq_528 <= _greatereq_data_528;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1925__delay_1924__variable_512 <= __delay_data_1924__variable_512;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1928__delay_1927__variable_513 <= __delay_data_1927__variable_513;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1931__delay_1930__variable_514 <= __delay_data_1930__variable_514;
      end 
      if(_mul_24_stream_oready) begin
        _cond_data_525 <= (__delay_data_1921_greaterthan_515)? _sll_data_519 : 1'sd0;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1923__delay_1922_greatereq_528 <= __delay_data_1922_greatereq_528;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1926__delay_1925__delay_1924__variable_512 <= __delay_data_1925__delay_1924__variable_512;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1929__delay_1928__delay_1927__variable_513 <= __delay_data_1928__delay_1927__variable_513;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1932__delay_1931__delay_1930__variable_514 <= __delay_data_1931__delay_1930__variable_514;
      end 
      if(_mul_24_stream_oready) begin
        __muladd_madd_odata_reg_531 <= __muladd_madd_odata_531;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1933__delay_1932__delay_1931____variable_514 <= __delay_data_1932__delay_1931__delay_1930__variable_514;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1934__delay_1933__delay_1932____variable_514 <= __delay_data_1933__delay_1932__delay_1931____variable_514;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1935__delay_1934__delay_1933____variable_514 <= __delay_data_1934__delay_1933__delay_1932____variable_514;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_1936__delay_1935__delay_1934____variable_514 <= __delay_data_1935__delay_1934__delay_1933____variable_514;
      end 
      if(_mul_24_stream_oready) begin
        _sra_data_532 <= __muladd_data_531 >>> __delay_data_1936__delay_1935__delay_1934____variable_514;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_512 <= _cond_data_1784;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_513 <= _cond_data_1451;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_514 <= __delay_data_2790__delay_2789_plus_1937;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1032 <= _mul_24_source_start;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1033 <= _tmp_1032;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1034 <= _tmp_1033;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1035 <= _mul_24_source_start;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1036 <= _tmp_1035;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1037 <= _tmp_1036;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1038 <= _tmp_1037;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1039 <= _tmp_1038;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1040 <= _tmp_1039;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1041 <= _tmp_1040;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1042 <= _tmp_1041;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1043 <= _tmp_1042;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1044 <= _tmp_1043;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1045 <= _mul_24_source_stop;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1046 <= _tmp_1045;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1047 <= _tmp_1046;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1048 <= _tmp_1047;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1049 <= _tmp_1048;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1050 <= _tmp_1049;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1051 <= _tmp_1050;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1052 <= _tmp_1051;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1053 <= _tmp_1052;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1054 <= _tmp_1053;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1055 <= _mul_24_source_busy;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1056 <= _tmp_1055;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1057 <= _tmp_1056;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1058 <= _tmp_1057;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1059 <= _tmp_1058;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1060 <= _tmp_1059;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1061 <= _tmp_1060;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1062 <= _tmp_1061;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1063 <= _tmp_1062;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1064 <= _tmp_1063;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_1065 <= _mul_24_sink_busy;
      end 
      if(!_mul_24_sink_busy && _tmp_1065) begin
        _mul_24_busy_reg <= 0;
      end 
      if(_mul_24_source_busy) begin
        _mul_24_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_24_fsm_1 = 1;
  localparam _mul_24_fsm_2 = 2;
  localparam _mul_24_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_24_fsm <= _mul_24_fsm_init;
      _mul_24_source_start <= 0;
      _mul_24_source_busy <= 0;
      _mul_24_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_24_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_24_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_24_stream_oready && _tmp_1034) begin
        _mul_24_stream_ivalid <= 1;
      end 
      if(_mul_24_stream_oready && 1'd0) begin
        _mul_24_stream_ivalid <= 0;
      end 
      case(_mul_24_fsm)
        _mul_24_fsm_init: begin
          if(_mul_24_run_flag) begin
            _mul_24_source_start <= 1;
          end 
          if(_mul_24_run_flag) begin
            _mul_24_fsm <= _mul_24_fsm_1;
          end 
        end
        _mul_24_fsm_1: begin
          if(_mul_24_source_start && _mul_24_stream_oready) begin
            _mul_24_source_start <= 0;
            _mul_24_source_busy <= 1;
          end 
          if(_mul_24_source_start && _mul_24_stream_oready) begin
            _mul_24_fsm <= _mul_24_fsm_2;
          end 
        end
        _mul_24_fsm_2: begin
          if(_mul_24_stream_oready) begin
            _mul_24_fsm <= _mul_24_fsm_3;
          end 
        end
        _mul_24_fsm_3: begin
          if(_mul_24_stream_oready && 1'd0) begin
            _mul_24_source_busy <= 0;
          end 
          if(_mul_24_stream_oready && 1'd0 && _mul_24_run_flag) begin
            _mul_24_source_start <= 1;
          end 
          if(_mul_24_stream_oready && 1'd0) begin
            _mul_24_fsm <= _mul_24_fsm_init;
          end 
          if(_mul_24_stream_oready && 1'd0 && _mul_24_run_flag) begin
            _mul_24_fsm <= _mul_24_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_25_x_source_ram_renable <= 0;
      _mul_25_x_source_fifo_deq <= 0;
      _mul_25_x_idle <= 1;
      _mul_25_y_source_ram_renable <= 0;
      _mul_25_y_source_fifo_deq <= 0;
      _mul_25_y_idle <= 1;
      _mul_25_rshift_source_ram_renable <= 0;
      _mul_25_rshift_source_fifo_deq <= 0;
      _mul_25_rshift_idle <= 1;
      _mul_25_z_sink_wenable <= 0;
      _mul_25_z_sink_fifo_enq <= 0;
      __mul_25_stream_ivalid_1 <= 0;
      __mul_25_stream_ivalid_2 <= 0;
      __mul_25_stream_ivalid_3 <= 0;
      __mul_25_stream_ivalid_4 <= 0;
      __mul_25_stream_ivalid_5 <= 0;
      __mul_25_stream_ivalid_6 <= 0;
      __mul_25_stream_ivalid_7 <= 0;
      __mul_25_stream_ivalid_8 <= 0;
      _greaterthan_data_536 <= 0;
      _minus_data_538 <= 0;
      _greatereq_data_549 <= 0;
      __delay_data_1943__variable_533 <= 0;
      __delay_data_1946__variable_534 <= 0;
      __delay_data_1949__variable_535 <= 0;
      _sll_data_540 <= 0;
      __delay_data_1940_greaterthan_536 <= 0;
      __delay_data_1941_greatereq_549 <= 0;
      __delay_data_1944__delay_1943__variable_533 <= 0;
      __delay_data_1947__delay_1946__variable_534 <= 0;
      __delay_data_1950__delay_1949__variable_535 <= 0;
      _cond_data_546 <= 0;
      __delay_data_1942__delay_1941_greatereq_549 <= 0;
      __delay_data_1945__delay_1944__delay_1943__variable_533 <= 0;
      __delay_data_1948__delay_1947__delay_1946__variable_534 <= 0;
      __delay_data_1951__delay_1950__delay_1949__variable_535 <= 0;
      __muladd_madd_odata_reg_552 <= 0;
      __delay_data_1952__delay_1951__delay_1950____variable_535 <= 0;
      __delay_data_1953__delay_1952__delay_1951____variable_535 <= 0;
      __delay_data_1954__delay_1953__delay_1952____variable_535 <= 0;
      __delay_data_1955__delay_1954__delay_1953____variable_535 <= 0;
      _sra_data_553 <= 0;
      __variable_wdata_533 <= 0;
      __variable_wdata_534 <= 0;
      __variable_wdata_535 <= 0;
      _tmp_1066 <= 0;
      _tmp_1067 <= 0;
      _tmp_1068 <= 0;
      _tmp_1069 <= 0;
      _tmp_1070 <= 0;
      _tmp_1071 <= 0;
      _tmp_1072 <= 0;
      _tmp_1073 <= 0;
      _tmp_1074 <= 0;
      _tmp_1075 <= 0;
      _tmp_1076 <= 0;
      _tmp_1077 <= 0;
      _tmp_1078 <= 0;
      _tmp_1079 <= 0;
      _tmp_1080 <= 0;
      _tmp_1081 <= 0;
      _tmp_1082 <= 0;
      _tmp_1083 <= 0;
      _tmp_1084 <= 0;
      _tmp_1085 <= 0;
      _tmp_1086 <= 0;
      _tmp_1087 <= 0;
      _tmp_1088 <= 0;
      _tmp_1089 <= 0;
      _tmp_1090 <= 0;
      _tmp_1091 <= 0;
      _tmp_1092 <= 0;
      _tmp_1093 <= 0;
      _tmp_1094 <= 0;
      _tmp_1095 <= 0;
      _tmp_1096 <= 0;
      _tmp_1097 <= 0;
      _tmp_1098 <= 0;
      _tmp_1099 <= 0;
      _mul_25_busy_reg <= 0;
    end else begin
      if(_mul_25_stream_oready) begin
        _mul_25_x_source_ram_renable <= 0;
        _mul_25_x_source_fifo_deq <= 0;
      end 
      _mul_25_x_idle <= _mul_25_x_idle;
      if(_mul_25_stream_oready) begin
        _mul_25_y_source_ram_renable <= 0;
        _mul_25_y_source_fifo_deq <= 0;
      end 
      _mul_25_y_idle <= _mul_25_y_idle;
      if(_mul_25_stream_oready) begin
        _mul_25_rshift_source_ram_renable <= 0;
        _mul_25_rshift_source_fifo_deq <= 0;
      end 
      _mul_25_rshift_idle <= _mul_25_rshift_idle;
      if(_mul_25_stream_oready) begin
        _mul_25_z_sink_wenable <= 0;
        _mul_25_z_sink_fifo_enq <= 0;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_1 <= _mul_25_stream_ivalid;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_2 <= __mul_25_stream_ivalid_1;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_3 <= __mul_25_stream_ivalid_2;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_4 <= __mul_25_stream_ivalid_3;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_5 <= __mul_25_stream_ivalid_4;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_6 <= __mul_25_stream_ivalid_5;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_7 <= __mul_25_stream_ivalid_6;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_8 <= __mul_25_stream_ivalid_7;
      end 
      if(_mul_25_stream_oready) begin
        _greaterthan_data_536 <= mul_25_rshift_data > 1'sd0;
      end 
      if(_mul_25_stream_oready) begin
        _minus_data_538 <= mul_25_rshift_data - 2'sd1;
      end 
      if(_mul_25_stream_oready) begin
        _greatereq_data_549 <= mul_25_x_data >= 1'sd0;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1943__variable_533 <= mul_25_x_data;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1946__variable_534 <= mul_25_y_data;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1949__variable_535 <= mul_25_rshift_data;
      end 
      if(_mul_25_stream_oready) begin
        _sll_data_540 <= 2'sd1 << _minus_data_538;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1940_greaterthan_536 <= _greaterthan_data_536;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1941_greatereq_549 <= _greatereq_data_549;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1944__delay_1943__variable_533 <= __delay_data_1943__variable_533;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1947__delay_1946__variable_534 <= __delay_data_1946__variable_534;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1950__delay_1949__variable_535 <= __delay_data_1949__variable_535;
      end 
      if(_mul_25_stream_oready) begin
        _cond_data_546 <= (__delay_data_1940_greaterthan_536)? _sll_data_540 : 1'sd0;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1942__delay_1941_greatereq_549 <= __delay_data_1941_greatereq_549;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1945__delay_1944__delay_1943__variable_533 <= __delay_data_1944__delay_1943__variable_533;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1948__delay_1947__delay_1946__variable_534 <= __delay_data_1947__delay_1946__variable_534;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1951__delay_1950__delay_1949__variable_535 <= __delay_data_1950__delay_1949__variable_535;
      end 
      if(_mul_25_stream_oready) begin
        __muladd_madd_odata_reg_552 <= __muladd_madd_odata_552;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1952__delay_1951__delay_1950____variable_535 <= __delay_data_1951__delay_1950__delay_1949__variable_535;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1953__delay_1952__delay_1951____variable_535 <= __delay_data_1952__delay_1951__delay_1950____variable_535;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1954__delay_1953__delay_1952____variable_535 <= __delay_data_1953__delay_1952__delay_1951____variable_535;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_1955__delay_1954__delay_1953____variable_535 <= __delay_data_1954__delay_1953__delay_1952____variable_535;
      end 
      if(_mul_25_stream_oready) begin
        _sra_data_553 <= __muladd_data_552 >>> __delay_data_1955__delay_1954__delay_1953____variable_535;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_533 <= _cond_data_1786;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_534 <= _cond_data_1453;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_535 <= __delay_data_2807__delay_2806_plus_1956;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1066 <= _mul_25_source_start;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1067 <= _tmp_1066;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1068 <= _tmp_1067;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1069 <= _mul_25_source_start;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1070 <= _tmp_1069;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1071 <= _tmp_1070;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1072 <= _tmp_1071;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1073 <= _tmp_1072;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1074 <= _tmp_1073;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1075 <= _tmp_1074;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1076 <= _tmp_1075;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1077 <= _tmp_1076;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1078 <= _tmp_1077;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1079 <= _mul_25_source_stop;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1080 <= _tmp_1079;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1081 <= _tmp_1080;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1082 <= _tmp_1081;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1083 <= _tmp_1082;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1084 <= _tmp_1083;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1085 <= _tmp_1084;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1086 <= _tmp_1085;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1087 <= _tmp_1086;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1088 <= _tmp_1087;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1089 <= _mul_25_source_busy;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1090 <= _tmp_1089;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1091 <= _tmp_1090;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1092 <= _tmp_1091;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1093 <= _tmp_1092;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1094 <= _tmp_1093;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1095 <= _tmp_1094;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1096 <= _tmp_1095;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1097 <= _tmp_1096;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1098 <= _tmp_1097;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_1099 <= _mul_25_sink_busy;
      end 
      if(!_mul_25_sink_busy && _tmp_1099) begin
        _mul_25_busy_reg <= 0;
      end 
      if(_mul_25_source_busy) begin
        _mul_25_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_25_fsm_1 = 1;
  localparam _mul_25_fsm_2 = 2;
  localparam _mul_25_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_25_fsm <= _mul_25_fsm_init;
      _mul_25_source_start <= 0;
      _mul_25_source_busy <= 0;
      _mul_25_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_25_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_25_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_25_stream_oready && _tmp_1068) begin
        _mul_25_stream_ivalid <= 1;
      end 
      if(_mul_25_stream_oready && 1'd0) begin
        _mul_25_stream_ivalid <= 0;
      end 
      case(_mul_25_fsm)
        _mul_25_fsm_init: begin
          if(_mul_25_run_flag) begin
            _mul_25_source_start <= 1;
          end 
          if(_mul_25_run_flag) begin
            _mul_25_fsm <= _mul_25_fsm_1;
          end 
        end
        _mul_25_fsm_1: begin
          if(_mul_25_source_start && _mul_25_stream_oready) begin
            _mul_25_source_start <= 0;
            _mul_25_source_busy <= 1;
          end 
          if(_mul_25_source_start && _mul_25_stream_oready) begin
            _mul_25_fsm <= _mul_25_fsm_2;
          end 
        end
        _mul_25_fsm_2: begin
          if(_mul_25_stream_oready) begin
            _mul_25_fsm <= _mul_25_fsm_3;
          end 
        end
        _mul_25_fsm_3: begin
          if(_mul_25_stream_oready && 1'd0) begin
            _mul_25_source_busy <= 0;
          end 
          if(_mul_25_stream_oready && 1'd0 && _mul_25_run_flag) begin
            _mul_25_source_start <= 1;
          end 
          if(_mul_25_stream_oready && 1'd0) begin
            _mul_25_fsm <= _mul_25_fsm_init;
          end 
          if(_mul_25_stream_oready && 1'd0 && _mul_25_run_flag) begin
            _mul_25_fsm <= _mul_25_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_26_x_source_ram_renable <= 0;
      _mul_26_x_source_fifo_deq <= 0;
      _mul_26_x_idle <= 1;
      _mul_26_y_source_ram_renable <= 0;
      _mul_26_y_source_fifo_deq <= 0;
      _mul_26_y_idle <= 1;
      _mul_26_rshift_source_ram_renable <= 0;
      _mul_26_rshift_source_fifo_deq <= 0;
      _mul_26_rshift_idle <= 1;
      _mul_26_z_sink_wenable <= 0;
      _mul_26_z_sink_fifo_enq <= 0;
      __mul_26_stream_ivalid_1 <= 0;
      __mul_26_stream_ivalid_2 <= 0;
      __mul_26_stream_ivalid_3 <= 0;
      __mul_26_stream_ivalid_4 <= 0;
      __mul_26_stream_ivalid_5 <= 0;
      __mul_26_stream_ivalid_6 <= 0;
      __mul_26_stream_ivalid_7 <= 0;
      __mul_26_stream_ivalid_8 <= 0;
      _greaterthan_data_557 <= 0;
      _minus_data_559 <= 0;
      _greatereq_data_570 <= 0;
      __delay_data_2020__variable_554 <= 0;
      __delay_data_2023__variable_555 <= 0;
      __delay_data_2026__variable_556 <= 0;
      _sll_data_561 <= 0;
      __delay_data_2017_greaterthan_557 <= 0;
      __delay_data_2018_greatereq_570 <= 0;
      __delay_data_2021__delay_2020__variable_554 <= 0;
      __delay_data_2024__delay_2023__variable_555 <= 0;
      __delay_data_2027__delay_2026__variable_556 <= 0;
      _cond_data_567 <= 0;
      __delay_data_2019__delay_2018_greatereq_570 <= 0;
      __delay_data_2022__delay_2021__delay_2020__variable_554 <= 0;
      __delay_data_2025__delay_2024__delay_2023__variable_555 <= 0;
      __delay_data_2028__delay_2027__delay_2026__variable_556 <= 0;
      __muladd_madd_odata_reg_573 <= 0;
      __delay_data_2029__delay_2028__delay_2027____variable_556 <= 0;
      __delay_data_2030__delay_2029__delay_2028____variable_556 <= 0;
      __delay_data_2031__delay_2030__delay_2029____variable_556 <= 0;
      __delay_data_2032__delay_2031__delay_2030____variable_556 <= 0;
      _sra_data_574 <= 0;
      __variable_wdata_554 <= 0;
      __variable_wdata_555 <= 0;
      __variable_wdata_556 <= 0;
      _tmp_1185 <= 0;
      _tmp_1186 <= 0;
      _tmp_1187 <= 0;
      _tmp_1188 <= 0;
      _tmp_1189 <= 0;
      _tmp_1190 <= 0;
      _tmp_1191 <= 0;
      _tmp_1192 <= 0;
      _tmp_1193 <= 0;
      _tmp_1194 <= 0;
      _tmp_1195 <= 0;
      _tmp_1196 <= 0;
      _tmp_1197 <= 0;
      _tmp_1198 <= 0;
      _tmp_1199 <= 0;
      _tmp_1200 <= 0;
      _tmp_1201 <= 0;
      _tmp_1202 <= 0;
      _tmp_1203 <= 0;
      _tmp_1204 <= 0;
      _tmp_1205 <= 0;
      _tmp_1206 <= 0;
      _tmp_1207 <= 0;
      _tmp_1208 <= 0;
      _tmp_1209 <= 0;
      _tmp_1210 <= 0;
      _tmp_1211 <= 0;
      _tmp_1212 <= 0;
      _tmp_1213 <= 0;
      _tmp_1214 <= 0;
      _tmp_1215 <= 0;
      _tmp_1216 <= 0;
      _tmp_1217 <= 0;
      _tmp_1218 <= 0;
      _mul_26_busy_reg <= 0;
    end else begin
      if(_mul_26_stream_oready) begin
        _mul_26_x_source_ram_renable <= 0;
        _mul_26_x_source_fifo_deq <= 0;
      end 
      _mul_26_x_idle <= _mul_26_x_idle;
      if(_mul_26_stream_oready) begin
        _mul_26_y_source_ram_renable <= 0;
        _mul_26_y_source_fifo_deq <= 0;
      end 
      _mul_26_y_idle <= _mul_26_y_idle;
      if(_mul_26_stream_oready) begin
        _mul_26_rshift_source_ram_renable <= 0;
        _mul_26_rshift_source_fifo_deq <= 0;
      end 
      _mul_26_rshift_idle <= _mul_26_rshift_idle;
      if(_mul_26_stream_oready) begin
        _mul_26_z_sink_wenable <= 0;
        _mul_26_z_sink_fifo_enq <= 0;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_1 <= _mul_26_stream_ivalid;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_2 <= __mul_26_stream_ivalid_1;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_3 <= __mul_26_stream_ivalid_2;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_4 <= __mul_26_stream_ivalid_3;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_5 <= __mul_26_stream_ivalid_4;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_6 <= __mul_26_stream_ivalid_5;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_7 <= __mul_26_stream_ivalid_6;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_8 <= __mul_26_stream_ivalid_7;
      end 
      if(_mul_26_stream_oready) begin
        _greaterthan_data_557 <= mul_26_rshift_data > 1'sd0;
      end 
      if(_mul_26_stream_oready) begin
        _minus_data_559 <= mul_26_rshift_data - 2'sd1;
      end 
      if(_mul_26_stream_oready) begin
        _greatereq_data_570 <= mul_26_x_data >= 1'sd0;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2020__variable_554 <= mul_26_x_data;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2023__variable_555 <= mul_26_y_data;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2026__variable_556 <= mul_26_rshift_data;
      end 
      if(_mul_26_stream_oready) begin
        _sll_data_561 <= 2'sd1 << _minus_data_559;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2017_greaterthan_557 <= _greaterthan_data_557;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2018_greatereq_570 <= _greatereq_data_570;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2021__delay_2020__variable_554 <= __delay_data_2020__variable_554;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2024__delay_2023__variable_555 <= __delay_data_2023__variable_555;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2027__delay_2026__variable_556 <= __delay_data_2026__variable_556;
      end 
      if(_mul_26_stream_oready) begin
        _cond_data_567 <= (__delay_data_2017_greaterthan_557)? _sll_data_561 : 1'sd0;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2019__delay_2018_greatereq_570 <= __delay_data_2018_greatereq_570;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2022__delay_2021__delay_2020__variable_554 <= __delay_data_2021__delay_2020__variable_554;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2025__delay_2024__delay_2023__variable_555 <= __delay_data_2024__delay_2023__variable_555;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2028__delay_2027__delay_2026__variable_556 <= __delay_data_2027__delay_2026__variable_556;
      end 
      if(_mul_26_stream_oready) begin
        __muladd_madd_odata_reg_573 <= __muladd_madd_odata_573;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2029__delay_2028__delay_2027____variable_556 <= __delay_data_2028__delay_2027__delay_2026__variable_556;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2030__delay_2029__delay_2028____variable_556 <= __delay_data_2029__delay_2028__delay_2027____variable_556;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2031__delay_2030__delay_2029____variable_556 <= __delay_data_2030__delay_2029__delay_2028____variable_556;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2032__delay_2031__delay_2030____variable_556 <= __delay_data_2031__delay_2030__delay_2029____variable_556;
      end 
      if(_mul_26_stream_oready) begin
        _sra_data_574 <= __muladd_data_573 >>> __delay_data_2032__delay_2031__delay_2030____variable_556;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_554 <= _cond_data_1999;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_555 <= _cond_data_1527;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_556 <= __delay_data_2859__delay_2858_plus_2033;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1185 <= _mul_26_source_start;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1186 <= _tmp_1185;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1187 <= _tmp_1186;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1188 <= _mul_26_source_start;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1189 <= _tmp_1188;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1190 <= _tmp_1189;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1191 <= _tmp_1190;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1192 <= _tmp_1191;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1193 <= _tmp_1192;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1194 <= _tmp_1193;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1195 <= _tmp_1194;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1196 <= _tmp_1195;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1197 <= _tmp_1196;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1198 <= _mul_26_source_stop;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1199 <= _tmp_1198;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1200 <= _tmp_1199;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1201 <= _tmp_1200;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1202 <= _tmp_1201;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1203 <= _tmp_1202;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1204 <= _tmp_1203;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1205 <= _tmp_1204;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1206 <= _tmp_1205;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1207 <= _tmp_1206;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1208 <= _mul_26_source_busy;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1209 <= _tmp_1208;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1210 <= _tmp_1209;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1211 <= _tmp_1210;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1212 <= _tmp_1211;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1213 <= _tmp_1212;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1214 <= _tmp_1213;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1215 <= _tmp_1214;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1216 <= _tmp_1215;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1217 <= _tmp_1216;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_1218 <= _mul_26_sink_busy;
      end 
      if(!_mul_26_sink_busy && _tmp_1218) begin
        _mul_26_busy_reg <= 0;
      end 
      if(_mul_26_source_busy) begin
        _mul_26_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_26_fsm_1 = 1;
  localparam _mul_26_fsm_2 = 2;
  localparam _mul_26_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_26_fsm <= _mul_26_fsm_init;
      _mul_26_source_start <= 0;
      _mul_26_source_busy <= 0;
      _mul_26_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_26_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_26_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_26_stream_oready && _tmp_1187) begin
        _mul_26_stream_ivalid <= 1;
      end 
      if(_mul_26_stream_oready && 1'd0) begin
        _mul_26_stream_ivalid <= 0;
      end 
      case(_mul_26_fsm)
        _mul_26_fsm_init: begin
          if(_mul_26_run_flag) begin
            _mul_26_source_start <= 1;
          end 
          if(_mul_26_run_flag) begin
            _mul_26_fsm <= _mul_26_fsm_1;
          end 
        end
        _mul_26_fsm_1: begin
          if(_mul_26_source_start && _mul_26_stream_oready) begin
            _mul_26_source_start <= 0;
            _mul_26_source_busy <= 1;
          end 
          if(_mul_26_source_start && _mul_26_stream_oready) begin
            _mul_26_fsm <= _mul_26_fsm_2;
          end 
        end
        _mul_26_fsm_2: begin
          if(_mul_26_stream_oready) begin
            _mul_26_fsm <= _mul_26_fsm_3;
          end 
        end
        _mul_26_fsm_3: begin
          if(_mul_26_stream_oready && 1'd0) begin
            _mul_26_source_busy <= 0;
          end 
          if(_mul_26_stream_oready && 1'd0 && _mul_26_run_flag) begin
            _mul_26_source_start <= 1;
          end 
          if(_mul_26_stream_oready && 1'd0) begin
            _mul_26_fsm <= _mul_26_fsm_init;
          end 
          if(_mul_26_stream_oready && 1'd0 && _mul_26_run_flag) begin
            _mul_26_fsm <= _mul_26_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_27_x_source_ram_renable <= 0;
      _mul_27_x_source_fifo_deq <= 0;
      _mul_27_x_idle <= 1;
      _mul_27_y_source_ram_renable <= 0;
      _mul_27_y_source_fifo_deq <= 0;
      _mul_27_y_idle <= 1;
      _mul_27_rshift_source_ram_renable <= 0;
      _mul_27_rshift_source_fifo_deq <= 0;
      _mul_27_rshift_idle <= 1;
      _mul_27_z_sink_wenable <= 0;
      _mul_27_z_sink_fifo_enq <= 0;
      __mul_27_stream_ivalid_1 <= 0;
      __mul_27_stream_ivalid_2 <= 0;
      __mul_27_stream_ivalid_3 <= 0;
      __mul_27_stream_ivalid_4 <= 0;
      __mul_27_stream_ivalid_5 <= 0;
      __mul_27_stream_ivalid_6 <= 0;
      __mul_27_stream_ivalid_7 <= 0;
      __mul_27_stream_ivalid_8 <= 0;
      _greaterthan_data_578 <= 0;
      _minus_data_580 <= 0;
      _greatereq_data_591 <= 0;
      __delay_data_2039__variable_575 <= 0;
      __delay_data_2042__variable_576 <= 0;
      __delay_data_2045__variable_577 <= 0;
      _sll_data_582 <= 0;
      __delay_data_2036_greaterthan_578 <= 0;
      __delay_data_2037_greatereq_591 <= 0;
      __delay_data_2040__delay_2039__variable_575 <= 0;
      __delay_data_2043__delay_2042__variable_576 <= 0;
      __delay_data_2046__delay_2045__variable_577 <= 0;
      _cond_data_588 <= 0;
      __delay_data_2038__delay_2037_greatereq_591 <= 0;
      __delay_data_2041__delay_2040__delay_2039__variable_575 <= 0;
      __delay_data_2044__delay_2043__delay_2042__variable_576 <= 0;
      __delay_data_2047__delay_2046__delay_2045__variable_577 <= 0;
      __muladd_madd_odata_reg_594 <= 0;
      __delay_data_2048__delay_2047__delay_2046____variable_577 <= 0;
      __delay_data_2049__delay_2048__delay_2047____variable_577 <= 0;
      __delay_data_2050__delay_2049__delay_2048____variable_577 <= 0;
      __delay_data_2051__delay_2050__delay_2049____variable_577 <= 0;
      _sra_data_595 <= 0;
      __variable_wdata_575 <= 0;
      __variable_wdata_576 <= 0;
      __variable_wdata_577 <= 0;
      _tmp_1219 <= 0;
      _tmp_1220 <= 0;
      _tmp_1221 <= 0;
      _tmp_1222 <= 0;
      _tmp_1223 <= 0;
      _tmp_1224 <= 0;
      _tmp_1225 <= 0;
      _tmp_1226 <= 0;
      _tmp_1227 <= 0;
      _tmp_1228 <= 0;
      _tmp_1229 <= 0;
      _tmp_1230 <= 0;
      _tmp_1231 <= 0;
      _tmp_1232 <= 0;
      _tmp_1233 <= 0;
      _tmp_1234 <= 0;
      _tmp_1235 <= 0;
      _tmp_1236 <= 0;
      _tmp_1237 <= 0;
      _tmp_1238 <= 0;
      _tmp_1239 <= 0;
      _tmp_1240 <= 0;
      _tmp_1241 <= 0;
      _tmp_1242 <= 0;
      _tmp_1243 <= 0;
      _tmp_1244 <= 0;
      _tmp_1245 <= 0;
      _tmp_1246 <= 0;
      _tmp_1247 <= 0;
      _tmp_1248 <= 0;
      _tmp_1249 <= 0;
      _tmp_1250 <= 0;
      _tmp_1251 <= 0;
      _tmp_1252 <= 0;
      _mul_27_busy_reg <= 0;
    end else begin
      if(_mul_27_stream_oready) begin
        _mul_27_x_source_ram_renable <= 0;
        _mul_27_x_source_fifo_deq <= 0;
      end 
      _mul_27_x_idle <= _mul_27_x_idle;
      if(_mul_27_stream_oready) begin
        _mul_27_y_source_ram_renable <= 0;
        _mul_27_y_source_fifo_deq <= 0;
      end 
      _mul_27_y_idle <= _mul_27_y_idle;
      if(_mul_27_stream_oready) begin
        _mul_27_rshift_source_ram_renable <= 0;
        _mul_27_rshift_source_fifo_deq <= 0;
      end 
      _mul_27_rshift_idle <= _mul_27_rshift_idle;
      if(_mul_27_stream_oready) begin
        _mul_27_z_sink_wenable <= 0;
        _mul_27_z_sink_fifo_enq <= 0;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_1 <= _mul_27_stream_ivalid;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_2 <= __mul_27_stream_ivalid_1;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_3 <= __mul_27_stream_ivalid_2;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_4 <= __mul_27_stream_ivalid_3;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_5 <= __mul_27_stream_ivalid_4;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_6 <= __mul_27_stream_ivalid_5;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_7 <= __mul_27_stream_ivalid_6;
      end 
      if(_mul_27_stream_oready) begin
        __mul_27_stream_ivalid_8 <= __mul_27_stream_ivalid_7;
      end 
      if(_mul_27_stream_oready) begin
        _greaterthan_data_578 <= mul_27_rshift_data > 1'sd0;
      end 
      if(_mul_27_stream_oready) begin
        _minus_data_580 <= mul_27_rshift_data - 2'sd1;
      end 
      if(_mul_27_stream_oready) begin
        _greatereq_data_591 <= mul_27_x_data >= 1'sd0;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2039__variable_575 <= mul_27_x_data;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2042__variable_576 <= mul_27_y_data;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2045__variable_577 <= mul_27_rshift_data;
      end 
      if(_mul_27_stream_oready) begin
        _sll_data_582 <= 2'sd1 << _minus_data_580;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2036_greaterthan_578 <= _greaterthan_data_578;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2037_greatereq_591 <= _greatereq_data_591;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2040__delay_2039__variable_575 <= __delay_data_2039__variable_575;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2043__delay_2042__variable_576 <= __delay_data_2042__variable_576;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2046__delay_2045__variable_577 <= __delay_data_2045__variable_577;
      end 
      if(_mul_27_stream_oready) begin
        _cond_data_588 <= (__delay_data_2036_greaterthan_578)? _sll_data_582 : 1'sd0;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2038__delay_2037_greatereq_591 <= __delay_data_2037_greatereq_591;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2041__delay_2040__delay_2039__variable_575 <= __delay_data_2040__delay_2039__variable_575;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2044__delay_2043__delay_2042__variable_576 <= __delay_data_2043__delay_2042__variable_576;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2047__delay_2046__delay_2045__variable_577 <= __delay_data_2046__delay_2045__variable_577;
      end 
      if(_mul_27_stream_oready) begin
        __muladd_madd_odata_reg_594 <= __muladd_madd_odata_594;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2048__delay_2047__delay_2046____variable_577 <= __delay_data_2047__delay_2046__delay_2045__variable_577;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2049__delay_2048__delay_2047____variable_577 <= __delay_data_2048__delay_2047__delay_2046____variable_577;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2050__delay_2049__delay_2048____variable_577 <= __delay_data_2049__delay_2048__delay_2047____variable_577;
      end 
      if(_mul_27_stream_oready) begin
        __delay_data_2051__delay_2050__delay_2049____variable_577 <= __delay_data_2050__delay_2049__delay_2048____variable_577;
      end 
      if(_mul_27_stream_oready) begin
        _sra_data_595 <= __muladd_data_594 >>> __delay_data_2051__delay_2050__delay_2049____variable_577;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_575 <= _cond_data_2001;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_576 <= _cond_data_1529;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_577 <= __delay_data_2869__delay_2868_plus_2052;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1219 <= _mul_27_source_start;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1220 <= _tmp_1219;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1221 <= _tmp_1220;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1222 <= _mul_27_source_start;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1223 <= _tmp_1222;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1224 <= _tmp_1223;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1225 <= _tmp_1224;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1226 <= _tmp_1225;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1227 <= _tmp_1226;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1228 <= _tmp_1227;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1229 <= _tmp_1228;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1230 <= _tmp_1229;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1231 <= _tmp_1230;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1232 <= _mul_27_source_stop;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1233 <= _tmp_1232;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1234 <= _tmp_1233;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1235 <= _tmp_1234;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1236 <= _tmp_1235;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1237 <= _tmp_1236;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1238 <= _tmp_1237;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1239 <= _tmp_1238;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1240 <= _tmp_1239;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1241 <= _tmp_1240;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1242 <= _mul_27_source_busy;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1243 <= _tmp_1242;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1244 <= _tmp_1243;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1245 <= _tmp_1244;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1246 <= _tmp_1245;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1247 <= _tmp_1246;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1248 <= _tmp_1247;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1249 <= _tmp_1248;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1250 <= _tmp_1249;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1251 <= _tmp_1250;
      end 
      if(_mul_27_stream_oready) begin
        _tmp_1252 <= _mul_27_sink_busy;
      end 
      if(!_mul_27_sink_busy && _tmp_1252) begin
        _mul_27_busy_reg <= 0;
      end 
      if(_mul_27_source_busy) begin
        _mul_27_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_27_fsm_1 = 1;
  localparam _mul_27_fsm_2 = 2;
  localparam _mul_27_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_27_fsm <= _mul_27_fsm_init;
      _mul_27_source_start <= 0;
      _mul_27_source_busy <= 0;
      _mul_27_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_27_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_27_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_27_stream_oready && _tmp_1221) begin
        _mul_27_stream_ivalid <= 1;
      end 
      if(_mul_27_stream_oready && 1'd0) begin
        _mul_27_stream_ivalid <= 0;
      end 
      case(_mul_27_fsm)
        _mul_27_fsm_init: begin
          if(_mul_27_run_flag) begin
            _mul_27_source_start <= 1;
          end 
          if(_mul_27_run_flag) begin
            _mul_27_fsm <= _mul_27_fsm_1;
          end 
        end
        _mul_27_fsm_1: begin
          if(_mul_27_source_start && _mul_27_stream_oready) begin
            _mul_27_source_start <= 0;
            _mul_27_source_busy <= 1;
          end 
          if(_mul_27_source_start && _mul_27_stream_oready) begin
            _mul_27_fsm <= _mul_27_fsm_2;
          end 
        end
        _mul_27_fsm_2: begin
          if(_mul_27_stream_oready) begin
            _mul_27_fsm <= _mul_27_fsm_3;
          end 
        end
        _mul_27_fsm_3: begin
          if(_mul_27_stream_oready && 1'd0) begin
            _mul_27_source_busy <= 0;
          end 
          if(_mul_27_stream_oready && 1'd0 && _mul_27_run_flag) begin
            _mul_27_source_start <= 1;
          end 
          if(_mul_27_stream_oready && 1'd0) begin
            _mul_27_fsm <= _mul_27_fsm_init;
          end 
          if(_mul_27_stream_oready && 1'd0 && _mul_27_run_flag) begin
            _mul_27_fsm <= _mul_27_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_28_x_source_ram_renable <= 0;
      _mul_28_x_source_fifo_deq <= 0;
      _mul_28_x_idle <= 1;
      _mul_28_y_source_ram_renable <= 0;
      _mul_28_y_source_fifo_deq <= 0;
      _mul_28_y_idle <= 1;
      _mul_28_rshift_source_ram_renable <= 0;
      _mul_28_rshift_source_fifo_deq <= 0;
      _mul_28_rshift_idle <= 1;
      _mul_28_z_sink_wenable <= 0;
      _mul_28_z_sink_fifo_enq <= 0;
      __mul_28_stream_ivalid_1 <= 0;
      __mul_28_stream_ivalid_2 <= 0;
      __mul_28_stream_ivalid_3 <= 0;
      __mul_28_stream_ivalid_4 <= 0;
      __mul_28_stream_ivalid_5 <= 0;
      __mul_28_stream_ivalid_6 <= 0;
      __mul_28_stream_ivalid_7 <= 0;
      __mul_28_stream_ivalid_8 <= 0;
      _greaterthan_data_599 <= 0;
      _minus_data_601 <= 0;
      _greatereq_data_612 <= 0;
      __delay_data_2058__variable_596 <= 0;
      __delay_data_2061__variable_597 <= 0;
      __delay_data_2064__variable_598 <= 0;
      _sll_data_603 <= 0;
      __delay_data_2055_greaterthan_599 <= 0;
      __delay_data_2056_greatereq_612 <= 0;
      __delay_data_2059__delay_2058__variable_596 <= 0;
      __delay_data_2062__delay_2061__variable_597 <= 0;
      __delay_data_2065__delay_2064__variable_598 <= 0;
      _cond_data_609 <= 0;
      __delay_data_2057__delay_2056_greatereq_612 <= 0;
      __delay_data_2060__delay_2059__delay_2058__variable_596 <= 0;
      __delay_data_2063__delay_2062__delay_2061__variable_597 <= 0;
      __delay_data_2066__delay_2065__delay_2064__variable_598 <= 0;
      __muladd_madd_odata_reg_615 <= 0;
      __delay_data_2067__delay_2066__delay_2065____variable_598 <= 0;
      __delay_data_2068__delay_2067__delay_2066____variable_598 <= 0;
      __delay_data_2069__delay_2068__delay_2067____variable_598 <= 0;
      __delay_data_2070__delay_2069__delay_2068____variable_598 <= 0;
      _sra_data_616 <= 0;
      __variable_wdata_596 <= 0;
      __variable_wdata_597 <= 0;
      __variable_wdata_598 <= 0;
      _tmp_1253 <= 0;
      _tmp_1254 <= 0;
      _tmp_1255 <= 0;
      _tmp_1256 <= 0;
      _tmp_1257 <= 0;
      _tmp_1258 <= 0;
      _tmp_1259 <= 0;
      _tmp_1260 <= 0;
      _tmp_1261 <= 0;
      _tmp_1262 <= 0;
      _tmp_1263 <= 0;
      _tmp_1264 <= 0;
      _tmp_1265 <= 0;
      _tmp_1266 <= 0;
      _tmp_1267 <= 0;
      _tmp_1268 <= 0;
      _tmp_1269 <= 0;
      _tmp_1270 <= 0;
      _tmp_1271 <= 0;
      _tmp_1272 <= 0;
      _tmp_1273 <= 0;
      _tmp_1274 <= 0;
      _tmp_1275 <= 0;
      _tmp_1276 <= 0;
      _tmp_1277 <= 0;
      _tmp_1278 <= 0;
      _tmp_1279 <= 0;
      _tmp_1280 <= 0;
      _tmp_1281 <= 0;
      _tmp_1282 <= 0;
      _tmp_1283 <= 0;
      _tmp_1284 <= 0;
      _tmp_1285 <= 0;
      _tmp_1286 <= 0;
      _mul_28_busy_reg <= 0;
    end else begin
      if(_mul_28_stream_oready) begin
        _mul_28_x_source_ram_renable <= 0;
        _mul_28_x_source_fifo_deq <= 0;
      end 
      _mul_28_x_idle <= _mul_28_x_idle;
      if(_mul_28_stream_oready) begin
        _mul_28_y_source_ram_renable <= 0;
        _mul_28_y_source_fifo_deq <= 0;
      end 
      _mul_28_y_idle <= _mul_28_y_idle;
      if(_mul_28_stream_oready) begin
        _mul_28_rshift_source_ram_renable <= 0;
        _mul_28_rshift_source_fifo_deq <= 0;
      end 
      _mul_28_rshift_idle <= _mul_28_rshift_idle;
      if(_mul_28_stream_oready) begin
        _mul_28_z_sink_wenable <= 0;
        _mul_28_z_sink_fifo_enq <= 0;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_1 <= _mul_28_stream_ivalid;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_2 <= __mul_28_stream_ivalid_1;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_3 <= __mul_28_stream_ivalid_2;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_4 <= __mul_28_stream_ivalid_3;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_5 <= __mul_28_stream_ivalid_4;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_6 <= __mul_28_stream_ivalid_5;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_7 <= __mul_28_stream_ivalid_6;
      end 
      if(_mul_28_stream_oready) begin
        __mul_28_stream_ivalid_8 <= __mul_28_stream_ivalid_7;
      end 
      if(_mul_28_stream_oready) begin
        _greaterthan_data_599 <= mul_28_rshift_data > 1'sd0;
      end 
      if(_mul_28_stream_oready) begin
        _minus_data_601 <= mul_28_rshift_data - 2'sd1;
      end 
      if(_mul_28_stream_oready) begin
        _greatereq_data_612 <= mul_28_x_data >= 1'sd0;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2058__variable_596 <= mul_28_x_data;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2061__variable_597 <= mul_28_y_data;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2064__variable_598 <= mul_28_rshift_data;
      end 
      if(_mul_28_stream_oready) begin
        _sll_data_603 <= 2'sd1 << _minus_data_601;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2055_greaterthan_599 <= _greaterthan_data_599;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2056_greatereq_612 <= _greatereq_data_612;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2059__delay_2058__variable_596 <= __delay_data_2058__variable_596;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2062__delay_2061__variable_597 <= __delay_data_2061__variable_597;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2065__delay_2064__variable_598 <= __delay_data_2064__variable_598;
      end 
      if(_mul_28_stream_oready) begin
        _cond_data_609 <= (__delay_data_2055_greaterthan_599)? _sll_data_603 : 1'sd0;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2057__delay_2056_greatereq_612 <= __delay_data_2056_greatereq_612;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2060__delay_2059__delay_2058__variable_596 <= __delay_data_2059__delay_2058__variable_596;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2063__delay_2062__delay_2061__variable_597 <= __delay_data_2062__delay_2061__variable_597;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2066__delay_2065__delay_2064__variable_598 <= __delay_data_2065__delay_2064__variable_598;
      end 
      if(_mul_28_stream_oready) begin
        __muladd_madd_odata_reg_615 <= __muladd_madd_odata_615;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2067__delay_2066__delay_2065____variable_598 <= __delay_data_2066__delay_2065__delay_2064__variable_598;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2068__delay_2067__delay_2066____variable_598 <= __delay_data_2067__delay_2066__delay_2065____variable_598;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2069__delay_2068__delay_2067____variable_598 <= __delay_data_2068__delay_2067__delay_2066____variable_598;
      end 
      if(_mul_28_stream_oready) begin
        __delay_data_2070__delay_2069__delay_2068____variable_598 <= __delay_data_2069__delay_2068__delay_2067____variable_598;
      end 
      if(_mul_28_stream_oready) begin
        _sra_data_616 <= __muladd_data_615 >>> __delay_data_2070__delay_2069__delay_2068____variable_598;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_596 <= _cond_data_2003;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_597 <= _cond_data_1531;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_598 <= __delay_data_2879__delay_2878_plus_2071;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1253 <= _mul_28_source_start;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1254 <= _tmp_1253;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1255 <= _tmp_1254;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1256 <= _mul_28_source_start;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1257 <= _tmp_1256;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1258 <= _tmp_1257;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1259 <= _tmp_1258;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1260 <= _tmp_1259;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1261 <= _tmp_1260;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1262 <= _tmp_1261;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1263 <= _tmp_1262;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1264 <= _tmp_1263;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1265 <= _tmp_1264;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1266 <= _mul_28_source_stop;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1267 <= _tmp_1266;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1268 <= _tmp_1267;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1269 <= _tmp_1268;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1270 <= _tmp_1269;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1271 <= _tmp_1270;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1272 <= _tmp_1271;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1273 <= _tmp_1272;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1274 <= _tmp_1273;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1275 <= _tmp_1274;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1276 <= _mul_28_source_busy;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1277 <= _tmp_1276;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1278 <= _tmp_1277;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1279 <= _tmp_1278;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1280 <= _tmp_1279;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1281 <= _tmp_1280;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1282 <= _tmp_1281;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1283 <= _tmp_1282;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1284 <= _tmp_1283;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1285 <= _tmp_1284;
      end 
      if(_mul_28_stream_oready) begin
        _tmp_1286 <= _mul_28_sink_busy;
      end 
      if(!_mul_28_sink_busy && _tmp_1286) begin
        _mul_28_busy_reg <= 0;
      end 
      if(_mul_28_source_busy) begin
        _mul_28_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_28_fsm_1 = 1;
  localparam _mul_28_fsm_2 = 2;
  localparam _mul_28_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_28_fsm <= _mul_28_fsm_init;
      _mul_28_source_start <= 0;
      _mul_28_source_busy <= 0;
      _mul_28_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_28_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_28_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_28_stream_oready && _tmp_1255) begin
        _mul_28_stream_ivalid <= 1;
      end 
      if(_mul_28_stream_oready && 1'd0) begin
        _mul_28_stream_ivalid <= 0;
      end 
      case(_mul_28_fsm)
        _mul_28_fsm_init: begin
          if(_mul_28_run_flag) begin
            _mul_28_source_start <= 1;
          end 
          if(_mul_28_run_flag) begin
            _mul_28_fsm <= _mul_28_fsm_1;
          end 
        end
        _mul_28_fsm_1: begin
          if(_mul_28_source_start && _mul_28_stream_oready) begin
            _mul_28_source_start <= 0;
            _mul_28_source_busy <= 1;
          end 
          if(_mul_28_source_start && _mul_28_stream_oready) begin
            _mul_28_fsm <= _mul_28_fsm_2;
          end 
        end
        _mul_28_fsm_2: begin
          if(_mul_28_stream_oready) begin
            _mul_28_fsm <= _mul_28_fsm_3;
          end 
        end
        _mul_28_fsm_3: begin
          if(_mul_28_stream_oready && 1'd0) begin
            _mul_28_source_busy <= 0;
          end 
          if(_mul_28_stream_oready && 1'd0 && _mul_28_run_flag) begin
            _mul_28_source_start <= 1;
          end 
          if(_mul_28_stream_oready && 1'd0) begin
            _mul_28_fsm <= _mul_28_fsm_init;
          end 
          if(_mul_28_stream_oready && 1'd0 && _mul_28_run_flag) begin
            _mul_28_fsm <= _mul_28_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_29_x_source_ram_renable <= 0;
      _mul_29_x_source_fifo_deq <= 0;
      _mul_29_x_idle <= 1;
      _mul_29_y_source_ram_renable <= 0;
      _mul_29_y_source_fifo_deq <= 0;
      _mul_29_y_idle <= 1;
      _mul_29_rshift_source_ram_renable <= 0;
      _mul_29_rshift_source_fifo_deq <= 0;
      _mul_29_rshift_idle <= 1;
      _mul_29_z_sink_wenable <= 0;
      _mul_29_z_sink_fifo_enq <= 0;
      __mul_29_stream_ivalid_1 <= 0;
      __mul_29_stream_ivalid_2 <= 0;
      __mul_29_stream_ivalid_3 <= 0;
      __mul_29_stream_ivalid_4 <= 0;
      __mul_29_stream_ivalid_5 <= 0;
      __mul_29_stream_ivalid_6 <= 0;
      __mul_29_stream_ivalid_7 <= 0;
      __mul_29_stream_ivalid_8 <= 0;
      _greaterthan_data_620 <= 0;
      _minus_data_622 <= 0;
      _greatereq_data_633 <= 0;
      __delay_data_2077__variable_617 <= 0;
      __delay_data_2080__variable_618 <= 0;
      __delay_data_2083__variable_619 <= 0;
      _sll_data_624 <= 0;
      __delay_data_2074_greaterthan_620 <= 0;
      __delay_data_2075_greatereq_633 <= 0;
      __delay_data_2078__delay_2077__variable_617 <= 0;
      __delay_data_2081__delay_2080__variable_618 <= 0;
      __delay_data_2084__delay_2083__variable_619 <= 0;
      _cond_data_630 <= 0;
      __delay_data_2076__delay_2075_greatereq_633 <= 0;
      __delay_data_2079__delay_2078__delay_2077__variable_617 <= 0;
      __delay_data_2082__delay_2081__delay_2080__variable_618 <= 0;
      __delay_data_2085__delay_2084__delay_2083__variable_619 <= 0;
      __muladd_madd_odata_reg_636 <= 0;
      __delay_data_2086__delay_2085__delay_2084____variable_619 <= 0;
      __delay_data_2087__delay_2086__delay_2085____variable_619 <= 0;
      __delay_data_2088__delay_2087__delay_2086____variable_619 <= 0;
      __delay_data_2089__delay_2088__delay_2087____variable_619 <= 0;
      _sra_data_637 <= 0;
      __variable_wdata_617 <= 0;
      __variable_wdata_618 <= 0;
      __variable_wdata_619 <= 0;
      _tmp_1287 <= 0;
      _tmp_1288 <= 0;
      _tmp_1289 <= 0;
      _tmp_1290 <= 0;
      _tmp_1291 <= 0;
      _tmp_1292 <= 0;
      _tmp_1293 <= 0;
      _tmp_1294 <= 0;
      _tmp_1295 <= 0;
      _tmp_1296 <= 0;
      _tmp_1297 <= 0;
      _tmp_1298 <= 0;
      _tmp_1299 <= 0;
      _tmp_1300 <= 0;
      _tmp_1301 <= 0;
      _tmp_1302 <= 0;
      _tmp_1303 <= 0;
      _tmp_1304 <= 0;
      _tmp_1305 <= 0;
      _tmp_1306 <= 0;
      _tmp_1307 <= 0;
      _tmp_1308 <= 0;
      _tmp_1309 <= 0;
      _tmp_1310 <= 0;
      _tmp_1311 <= 0;
      _tmp_1312 <= 0;
      _tmp_1313 <= 0;
      _tmp_1314 <= 0;
      _tmp_1315 <= 0;
      _tmp_1316 <= 0;
      _tmp_1317 <= 0;
      _tmp_1318 <= 0;
      _tmp_1319 <= 0;
      _tmp_1320 <= 0;
      _mul_29_busy_reg <= 0;
    end else begin
      if(_mul_29_stream_oready) begin
        _mul_29_x_source_ram_renable <= 0;
        _mul_29_x_source_fifo_deq <= 0;
      end 
      _mul_29_x_idle <= _mul_29_x_idle;
      if(_mul_29_stream_oready) begin
        _mul_29_y_source_ram_renable <= 0;
        _mul_29_y_source_fifo_deq <= 0;
      end 
      _mul_29_y_idle <= _mul_29_y_idle;
      if(_mul_29_stream_oready) begin
        _mul_29_rshift_source_ram_renable <= 0;
        _mul_29_rshift_source_fifo_deq <= 0;
      end 
      _mul_29_rshift_idle <= _mul_29_rshift_idle;
      if(_mul_29_stream_oready) begin
        _mul_29_z_sink_wenable <= 0;
        _mul_29_z_sink_fifo_enq <= 0;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_1 <= _mul_29_stream_ivalid;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_2 <= __mul_29_stream_ivalid_1;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_3 <= __mul_29_stream_ivalid_2;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_4 <= __mul_29_stream_ivalid_3;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_5 <= __mul_29_stream_ivalid_4;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_6 <= __mul_29_stream_ivalid_5;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_7 <= __mul_29_stream_ivalid_6;
      end 
      if(_mul_29_stream_oready) begin
        __mul_29_stream_ivalid_8 <= __mul_29_stream_ivalid_7;
      end 
      if(_mul_29_stream_oready) begin
        _greaterthan_data_620 <= mul_29_rshift_data > 1'sd0;
      end 
      if(_mul_29_stream_oready) begin
        _minus_data_622 <= mul_29_rshift_data - 2'sd1;
      end 
      if(_mul_29_stream_oready) begin
        _greatereq_data_633 <= mul_29_x_data >= 1'sd0;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2077__variable_617 <= mul_29_x_data;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2080__variable_618 <= mul_29_y_data;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2083__variable_619 <= mul_29_rshift_data;
      end 
      if(_mul_29_stream_oready) begin
        _sll_data_624 <= 2'sd1 << _minus_data_622;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2074_greaterthan_620 <= _greaterthan_data_620;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2075_greatereq_633 <= _greatereq_data_633;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2078__delay_2077__variable_617 <= __delay_data_2077__variable_617;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2081__delay_2080__variable_618 <= __delay_data_2080__variable_618;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2084__delay_2083__variable_619 <= __delay_data_2083__variable_619;
      end 
      if(_mul_29_stream_oready) begin
        _cond_data_630 <= (__delay_data_2074_greaterthan_620)? _sll_data_624 : 1'sd0;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2076__delay_2075_greatereq_633 <= __delay_data_2075_greatereq_633;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2079__delay_2078__delay_2077__variable_617 <= __delay_data_2078__delay_2077__variable_617;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2082__delay_2081__delay_2080__variable_618 <= __delay_data_2081__delay_2080__variable_618;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2085__delay_2084__delay_2083__variable_619 <= __delay_data_2084__delay_2083__variable_619;
      end 
      if(_mul_29_stream_oready) begin
        __muladd_madd_odata_reg_636 <= __muladd_madd_odata_636;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2086__delay_2085__delay_2084____variable_619 <= __delay_data_2085__delay_2084__delay_2083__variable_619;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2087__delay_2086__delay_2085____variable_619 <= __delay_data_2086__delay_2085__delay_2084____variable_619;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2088__delay_2087__delay_2086____variable_619 <= __delay_data_2087__delay_2086__delay_2085____variable_619;
      end 
      if(_mul_29_stream_oready) begin
        __delay_data_2089__delay_2088__delay_2087____variable_619 <= __delay_data_2088__delay_2087__delay_2086____variable_619;
      end 
      if(_mul_29_stream_oready) begin
        _sra_data_637 <= __muladd_data_636 >>> __delay_data_2089__delay_2088__delay_2087____variable_619;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_617 <= _cond_data_2005;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_618 <= _cond_data_1533;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_619 <= __delay_data_2889__delay_2888_plus_2090;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1287 <= _mul_29_source_start;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1288 <= _tmp_1287;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1289 <= _tmp_1288;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1290 <= _mul_29_source_start;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1291 <= _tmp_1290;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1292 <= _tmp_1291;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1293 <= _tmp_1292;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1294 <= _tmp_1293;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1295 <= _tmp_1294;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1296 <= _tmp_1295;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1297 <= _tmp_1296;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1298 <= _tmp_1297;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1299 <= _tmp_1298;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1300 <= _mul_29_source_stop;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1301 <= _tmp_1300;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1302 <= _tmp_1301;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1303 <= _tmp_1302;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1304 <= _tmp_1303;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1305 <= _tmp_1304;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1306 <= _tmp_1305;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1307 <= _tmp_1306;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1308 <= _tmp_1307;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1309 <= _tmp_1308;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1310 <= _mul_29_source_busy;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1311 <= _tmp_1310;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1312 <= _tmp_1311;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1313 <= _tmp_1312;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1314 <= _tmp_1313;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1315 <= _tmp_1314;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1316 <= _tmp_1315;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1317 <= _tmp_1316;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1318 <= _tmp_1317;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1319 <= _tmp_1318;
      end 
      if(_mul_29_stream_oready) begin
        _tmp_1320 <= _mul_29_sink_busy;
      end 
      if(!_mul_29_sink_busy && _tmp_1320) begin
        _mul_29_busy_reg <= 0;
      end 
      if(_mul_29_source_busy) begin
        _mul_29_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_29_fsm_1 = 1;
  localparam _mul_29_fsm_2 = 2;
  localparam _mul_29_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_29_fsm <= _mul_29_fsm_init;
      _mul_29_source_start <= 0;
      _mul_29_source_busy <= 0;
      _mul_29_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_29_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_29_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_29_stream_oready && _tmp_1289) begin
        _mul_29_stream_ivalid <= 1;
      end 
      if(_mul_29_stream_oready && 1'd0) begin
        _mul_29_stream_ivalid <= 0;
      end 
      case(_mul_29_fsm)
        _mul_29_fsm_init: begin
          if(_mul_29_run_flag) begin
            _mul_29_source_start <= 1;
          end 
          if(_mul_29_run_flag) begin
            _mul_29_fsm <= _mul_29_fsm_1;
          end 
        end
        _mul_29_fsm_1: begin
          if(_mul_29_source_start && _mul_29_stream_oready) begin
            _mul_29_source_start <= 0;
            _mul_29_source_busy <= 1;
          end 
          if(_mul_29_source_start && _mul_29_stream_oready) begin
            _mul_29_fsm <= _mul_29_fsm_2;
          end 
        end
        _mul_29_fsm_2: begin
          if(_mul_29_stream_oready) begin
            _mul_29_fsm <= _mul_29_fsm_3;
          end 
        end
        _mul_29_fsm_3: begin
          if(_mul_29_stream_oready && 1'd0) begin
            _mul_29_source_busy <= 0;
          end 
          if(_mul_29_stream_oready && 1'd0 && _mul_29_run_flag) begin
            _mul_29_source_start <= 1;
          end 
          if(_mul_29_stream_oready && 1'd0) begin
            _mul_29_fsm <= _mul_29_fsm_init;
          end 
          if(_mul_29_stream_oready && 1'd0 && _mul_29_run_flag) begin
            _mul_29_fsm <= _mul_29_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_30_x_source_ram_renable <= 0;
      _mul_30_x_source_fifo_deq <= 0;
      _mul_30_x_idle <= 1;
      _mul_30_y_source_ram_renable <= 0;
      _mul_30_y_source_fifo_deq <= 0;
      _mul_30_y_idle <= 1;
      _mul_30_rshift_source_ram_renable <= 0;
      _mul_30_rshift_source_fifo_deq <= 0;
      _mul_30_rshift_idle <= 1;
      _mul_30_z_sink_wenable <= 0;
      _mul_30_z_sink_fifo_enq <= 0;
      __mul_30_stream_ivalid_1 <= 0;
      __mul_30_stream_ivalid_2 <= 0;
      __mul_30_stream_ivalid_3 <= 0;
      __mul_30_stream_ivalid_4 <= 0;
      __mul_30_stream_ivalid_5 <= 0;
      __mul_30_stream_ivalid_6 <= 0;
      __mul_30_stream_ivalid_7 <= 0;
      __mul_30_stream_ivalid_8 <= 0;
      _greaterthan_data_641 <= 0;
      _minus_data_643 <= 0;
      _greatereq_data_654 <= 0;
      __delay_data_2096__variable_638 <= 0;
      __delay_data_2099__variable_639 <= 0;
      __delay_data_2102__variable_640 <= 0;
      _sll_data_645 <= 0;
      __delay_data_2093_greaterthan_641 <= 0;
      __delay_data_2094_greatereq_654 <= 0;
      __delay_data_2097__delay_2096__variable_638 <= 0;
      __delay_data_2100__delay_2099__variable_639 <= 0;
      __delay_data_2103__delay_2102__variable_640 <= 0;
      _cond_data_651 <= 0;
      __delay_data_2095__delay_2094_greatereq_654 <= 0;
      __delay_data_2098__delay_2097__delay_2096__variable_638 <= 0;
      __delay_data_2101__delay_2100__delay_2099__variable_639 <= 0;
      __delay_data_2104__delay_2103__delay_2102__variable_640 <= 0;
      __muladd_madd_odata_reg_657 <= 0;
      __delay_data_2105__delay_2104__delay_2103____variable_640 <= 0;
      __delay_data_2106__delay_2105__delay_2104____variable_640 <= 0;
      __delay_data_2107__delay_2106__delay_2105____variable_640 <= 0;
      __delay_data_2108__delay_2107__delay_2106____variable_640 <= 0;
      _sra_data_658 <= 0;
      __variable_wdata_638 <= 0;
      __variable_wdata_639 <= 0;
      __variable_wdata_640 <= 0;
      _tmp_1321 <= 0;
      _tmp_1322 <= 0;
      _tmp_1323 <= 0;
      _tmp_1324 <= 0;
      _tmp_1325 <= 0;
      _tmp_1326 <= 0;
      _tmp_1327 <= 0;
      _tmp_1328 <= 0;
      _tmp_1329 <= 0;
      _tmp_1330 <= 0;
      _tmp_1331 <= 0;
      _tmp_1332 <= 0;
      _tmp_1333 <= 0;
      _tmp_1334 <= 0;
      _tmp_1335 <= 0;
      _tmp_1336 <= 0;
      _tmp_1337 <= 0;
      _tmp_1338 <= 0;
      _tmp_1339 <= 0;
      _tmp_1340 <= 0;
      _tmp_1341 <= 0;
      _tmp_1342 <= 0;
      _tmp_1343 <= 0;
      _tmp_1344 <= 0;
      _tmp_1345 <= 0;
      _tmp_1346 <= 0;
      _tmp_1347 <= 0;
      _tmp_1348 <= 0;
      _tmp_1349 <= 0;
      _tmp_1350 <= 0;
      _tmp_1351 <= 0;
      _tmp_1352 <= 0;
      _tmp_1353 <= 0;
      _tmp_1354 <= 0;
      _mul_30_busy_reg <= 0;
    end else begin
      if(_mul_30_stream_oready) begin
        _mul_30_x_source_ram_renable <= 0;
        _mul_30_x_source_fifo_deq <= 0;
      end 
      _mul_30_x_idle <= _mul_30_x_idle;
      if(_mul_30_stream_oready) begin
        _mul_30_y_source_ram_renable <= 0;
        _mul_30_y_source_fifo_deq <= 0;
      end 
      _mul_30_y_idle <= _mul_30_y_idle;
      if(_mul_30_stream_oready) begin
        _mul_30_rshift_source_ram_renable <= 0;
        _mul_30_rshift_source_fifo_deq <= 0;
      end 
      _mul_30_rshift_idle <= _mul_30_rshift_idle;
      if(_mul_30_stream_oready) begin
        _mul_30_z_sink_wenable <= 0;
        _mul_30_z_sink_fifo_enq <= 0;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_1 <= _mul_30_stream_ivalid;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_2 <= __mul_30_stream_ivalid_1;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_3 <= __mul_30_stream_ivalid_2;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_4 <= __mul_30_stream_ivalid_3;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_5 <= __mul_30_stream_ivalid_4;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_6 <= __mul_30_stream_ivalid_5;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_7 <= __mul_30_stream_ivalid_6;
      end 
      if(_mul_30_stream_oready) begin
        __mul_30_stream_ivalid_8 <= __mul_30_stream_ivalid_7;
      end 
      if(_mul_30_stream_oready) begin
        _greaterthan_data_641 <= mul_30_rshift_data > 1'sd0;
      end 
      if(_mul_30_stream_oready) begin
        _minus_data_643 <= mul_30_rshift_data - 2'sd1;
      end 
      if(_mul_30_stream_oready) begin
        _greatereq_data_654 <= mul_30_x_data >= 1'sd0;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2096__variable_638 <= mul_30_x_data;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2099__variable_639 <= mul_30_y_data;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2102__variable_640 <= mul_30_rshift_data;
      end 
      if(_mul_30_stream_oready) begin
        _sll_data_645 <= 2'sd1 << _minus_data_643;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2093_greaterthan_641 <= _greaterthan_data_641;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2094_greatereq_654 <= _greatereq_data_654;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2097__delay_2096__variable_638 <= __delay_data_2096__variable_638;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2100__delay_2099__variable_639 <= __delay_data_2099__variable_639;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2103__delay_2102__variable_640 <= __delay_data_2102__variable_640;
      end 
      if(_mul_30_stream_oready) begin
        _cond_data_651 <= (__delay_data_2093_greaterthan_641)? _sll_data_645 : 1'sd0;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2095__delay_2094_greatereq_654 <= __delay_data_2094_greatereq_654;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2098__delay_2097__delay_2096__variable_638 <= __delay_data_2097__delay_2096__variable_638;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2101__delay_2100__delay_2099__variable_639 <= __delay_data_2100__delay_2099__variable_639;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2104__delay_2103__delay_2102__variable_640 <= __delay_data_2103__delay_2102__variable_640;
      end 
      if(_mul_30_stream_oready) begin
        __muladd_madd_odata_reg_657 <= __muladd_madd_odata_657;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2105__delay_2104__delay_2103____variable_640 <= __delay_data_2104__delay_2103__delay_2102__variable_640;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2106__delay_2105__delay_2104____variable_640 <= __delay_data_2105__delay_2104__delay_2103____variable_640;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2107__delay_2106__delay_2105____variable_640 <= __delay_data_2106__delay_2105__delay_2104____variable_640;
      end 
      if(_mul_30_stream_oready) begin
        __delay_data_2108__delay_2107__delay_2106____variable_640 <= __delay_data_2107__delay_2106__delay_2105____variable_640;
      end 
      if(_mul_30_stream_oready) begin
        _sra_data_658 <= __muladd_data_657 >>> __delay_data_2108__delay_2107__delay_2106____variable_640;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_638 <= _cond_data_2007;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_639 <= _cond_data_1535;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_640 <= __delay_data_2899__delay_2898_plus_2109;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1321 <= _mul_30_source_start;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1322 <= _tmp_1321;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1323 <= _tmp_1322;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1324 <= _mul_30_source_start;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1325 <= _tmp_1324;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1326 <= _tmp_1325;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1327 <= _tmp_1326;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1328 <= _tmp_1327;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1329 <= _tmp_1328;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1330 <= _tmp_1329;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1331 <= _tmp_1330;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1332 <= _tmp_1331;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1333 <= _tmp_1332;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1334 <= _mul_30_source_stop;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1335 <= _tmp_1334;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1336 <= _tmp_1335;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1337 <= _tmp_1336;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1338 <= _tmp_1337;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1339 <= _tmp_1338;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1340 <= _tmp_1339;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1341 <= _tmp_1340;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1342 <= _tmp_1341;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1343 <= _tmp_1342;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1344 <= _mul_30_source_busy;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1345 <= _tmp_1344;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1346 <= _tmp_1345;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1347 <= _tmp_1346;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1348 <= _tmp_1347;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1349 <= _tmp_1348;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1350 <= _tmp_1349;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1351 <= _tmp_1350;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1352 <= _tmp_1351;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1353 <= _tmp_1352;
      end 
      if(_mul_30_stream_oready) begin
        _tmp_1354 <= _mul_30_sink_busy;
      end 
      if(!_mul_30_sink_busy && _tmp_1354) begin
        _mul_30_busy_reg <= 0;
      end 
      if(_mul_30_source_busy) begin
        _mul_30_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_30_fsm_1 = 1;
  localparam _mul_30_fsm_2 = 2;
  localparam _mul_30_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_30_fsm <= _mul_30_fsm_init;
      _mul_30_source_start <= 0;
      _mul_30_source_busy <= 0;
      _mul_30_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_30_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_30_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_30_stream_oready && _tmp_1323) begin
        _mul_30_stream_ivalid <= 1;
      end 
      if(_mul_30_stream_oready && 1'd0) begin
        _mul_30_stream_ivalid <= 0;
      end 
      case(_mul_30_fsm)
        _mul_30_fsm_init: begin
          if(_mul_30_run_flag) begin
            _mul_30_source_start <= 1;
          end 
          if(_mul_30_run_flag) begin
            _mul_30_fsm <= _mul_30_fsm_1;
          end 
        end
        _mul_30_fsm_1: begin
          if(_mul_30_source_start && _mul_30_stream_oready) begin
            _mul_30_source_start <= 0;
            _mul_30_source_busy <= 1;
          end 
          if(_mul_30_source_start && _mul_30_stream_oready) begin
            _mul_30_fsm <= _mul_30_fsm_2;
          end 
        end
        _mul_30_fsm_2: begin
          if(_mul_30_stream_oready) begin
            _mul_30_fsm <= _mul_30_fsm_3;
          end 
        end
        _mul_30_fsm_3: begin
          if(_mul_30_stream_oready && 1'd0) begin
            _mul_30_source_busy <= 0;
          end 
          if(_mul_30_stream_oready && 1'd0 && _mul_30_run_flag) begin
            _mul_30_source_start <= 1;
          end 
          if(_mul_30_stream_oready && 1'd0) begin
            _mul_30_fsm <= _mul_30_fsm_init;
          end 
          if(_mul_30_stream_oready && 1'd0 && _mul_30_run_flag) begin
            _mul_30_fsm <= _mul_30_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_31_x_source_ram_renable <= 0;
      _mul_31_x_source_fifo_deq <= 0;
      _mul_31_x_idle <= 1;
      _mul_31_y_source_ram_renable <= 0;
      _mul_31_y_source_fifo_deq <= 0;
      _mul_31_y_idle <= 1;
      _mul_31_rshift_source_ram_renable <= 0;
      _mul_31_rshift_source_fifo_deq <= 0;
      _mul_31_rshift_idle <= 1;
      _mul_31_z_sink_wenable <= 0;
      _mul_31_z_sink_fifo_enq <= 0;
      __mul_31_stream_ivalid_1 <= 0;
      __mul_31_stream_ivalid_2 <= 0;
      __mul_31_stream_ivalid_3 <= 0;
      __mul_31_stream_ivalid_4 <= 0;
      __mul_31_stream_ivalid_5 <= 0;
      __mul_31_stream_ivalid_6 <= 0;
      __mul_31_stream_ivalid_7 <= 0;
      __mul_31_stream_ivalid_8 <= 0;
      _greaterthan_data_662 <= 0;
      _minus_data_664 <= 0;
      _greatereq_data_675 <= 0;
      __delay_data_2115__variable_659 <= 0;
      __delay_data_2118__variable_660 <= 0;
      __delay_data_2121__variable_661 <= 0;
      _sll_data_666 <= 0;
      __delay_data_2112_greaterthan_662 <= 0;
      __delay_data_2113_greatereq_675 <= 0;
      __delay_data_2116__delay_2115__variable_659 <= 0;
      __delay_data_2119__delay_2118__variable_660 <= 0;
      __delay_data_2122__delay_2121__variable_661 <= 0;
      _cond_data_672 <= 0;
      __delay_data_2114__delay_2113_greatereq_675 <= 0;
      __delay_data_2117__delay_2116__delay_2115__variable_659 <= 0;
      __delay_data_2120__delay_2119__delay_2118__variable_660 <= 0;
      __delay_data_2123__delay_2122__delay_2121__variable_661 <= 0;
      __muladd_madd_odata_reg_678 <= 0;
      __delay_data_2124__delay_2123__delay_2122____variable_661 <= 0;
      __delay_data_2125__delay_2124__delay_2123____variable_661 <= 0;
      __delay_data_2126__delay_2125__delay_2124____variable_661 <= 0;
      __delay_data_2127__delay_2126__delay_2125____variable_661 <= 0;
      _sra_data_679 <= 0;
      __variable_wdata_659 <= 0;
      __variable_wdata_660 <= 0;
      __variable_wdata_661 <= 0;
      _tmp_1355 <= 0;
      _tmp_1356 <= 0;
      _tmp_1357 <= 0;
      _tmp_1358 <= 0;
      _tmp_1359 <= 0;
      _tmp_1360 <= 0;
      _tmp_1361 <= 0;
      _tmp_1362 <= 0;
      _tmp_1363 <= 0;
      _tmp_1364 <= 0;
      _tmp_1365 <= 0;
      _tmp_1366 <= 0;
      _tmp_1367 <= 0;
      _tmp_1368 <= 0;
      _tmp_1369 <= 0;
      _tmp_1370 <= 0;
      _tmp_1371 <= 0;
      _tmp_1372 <= 0;
      _tmp_1373 <= 0;
      _tmp_1374 <= 0;
      _tmp_1375 <= 0;
      _tmp_1376 <= 0;
      _tmp_1377 <= 0;
      _tmp_1378 <= 0;
      _tmp_1379 <= 0;
      _tmp_1380 <= 0;
      _tmp_1381 <= 0;
      _tmp_1382 <= 0;
      _tmp_1383 <= 0;
      _tmp_1384 <= 0;
      _tmp_1385 <= 0;
      _tmp_1386 <= 0;
      _tmp_1387 <= 0;
      _tmp_1388 <= 0;
      _mul_31_busy_reg <= 0;
    end else begin
      if(_mul_31_stream_oready) begin
        _mul_31_x_source_ram_renable <= 0;
        _mul_31_x_source_fifo_deq <= 0;
      end 
      _mul_31_x_idle <= _mul_31_x_idle;
      if(_mul_31_stream_oready) begin
        _mul_31_y_source_ram_renable <= 0;
        _mul_31_y_source_fifo_deq <= 0;
      end 
      _mul_31_y_idle <= _mul_31_y_idle;
      if(_mul_31_stream_oready) begin
        _mul_31_rshift_source_ram_renable <= 0;
        _mul_31_rshift_source_fifo_deq <= 0;
      end 
      _mul_31_rshift_idle <= _mul_31_rshift_idle;
      if(_mul_31_stream_oready) begin
        _mul_31_z_sink_wenable <= 0;
        _mul_31_z_sink_fifo_enq <= 0;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_1 <= _mul_31_stream_ivalid;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_2 <= __mul_31_stream_ivalid_1;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_3 <= __mul_31_stream_ivalid_2;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_4 <= __mul_31_stream_ivalid_3;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_5 <= __mul_31_stream_ivalid_4;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_6 <= __mul_31_stream_ivalid_5;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_7 <= __mul_31_stream_ivalid_6;
      end 
      if(_mul_31_stream_oready) begin
        __mul_31_stream_ivalid_8 <= __mul_31_stream_ivalid_7;
      end 
      if(_mul_31_stream_oready) begin
        _greaterthan_data_662 <= mul_31_rshift_data > 1'sd0;
      end 
      if(_mul_31_stream_oready) begin
        _minus_data_664 <= mul_31_rshift_data - 2'sd1;
      end 
      if(_mul_31_stream_oready) begin
        _greatereq_data_675 <= mul_31_x_data >= 1'sd0;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2115__variable_659 <= mul_31_x_data;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2118__variable_660 <= mul_31_y_data;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2121__variable_661 <= mul_31_rshift_data;
      end 
      if(_mul_31_stream_oready) begin
        _sll_data_666 <= 2'sd1 << _minus_data_664;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2112_greaterthan_662 <= _greaterthan_data_662;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2113_greatereq_675 <= _greatereq_data_675;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2116__delay_2115__variable_659 <= __delay_data_2115__variable_659;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2119__delay_2118__variable_660 <= __delay_data_2118__variable_660;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2122__delay_2121__variable_661 <= __delay_data_2121__variable_661;
      end 
      if(_mul_31_stream_oready) begin
        _cond_data_672 <= (__delay_data_2112_greaterthan_662)? _sll_data_666 : 1'sd0;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2114__delay_2113_greatereq_675 <= __delay_data_2113_greatereq_675;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2117__delay_2116__delay_2115__variable_659 <= __delay_data_2116__delay_2115__variable_659;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2120__delay_2119__delay_2118__variable_660 <= __delay_data_2119__delay_2118__variable_660;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2123__delay_2122__delay_2121__variable_661 <= __delay_data_2122__delay_2121__variable_661;
      end 
      if(_mul_31_stream_oready) begin
        __muladd_madd_odata_reg_678 <= __muladd_madd_odata_678;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2124__delay_2123__delay_2122____variable_661 <= __delay_data_2123__delay_2122__delay_2121__variable_661;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2125__delay_2124__delay_2123____variable_661 <= __delay_data_2124__delay_2123__delay_2122____variable_661;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2126__delay_2125__delay_2124____variable_661 <= __delay_data_2125__delay_2124__delay_2123____variable_661;
      end 
      if(_mul_31_stream_oready) begin
        __delay_data_2127__delay_2126__delay_2125____variable_661 <= __delay_data_2126__delay_2125__delay_2124____variable_661;
      end 
      if(_mul_31_stream_oready) begin
        _sra_data_679 <= __muladd_data_678 >>> __delay_data_2127__delay_2126__delay_2125____variable_661;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_659 <= _cond_data_2009;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_660 <= _cond_data_1537;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_661 <= __delay_data_2909__delay_2908_plus_2128;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1355 <= _mul_31_source_start;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1356 <= _tmp_1355;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1357 <= _tmp_1356;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1358 <= _mul_31_source_start;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1359 <= _tmp_1358;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1360 <= _tmp_1359;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1361 <= _tmp_1360;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1362 <= _tmp_1361;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1363 <= _tmp_1362;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1364 <= _tmp_1363;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1365 <= _tmp_1364;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1366 <= _tmp_1365;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1367 <= _tmp_1366;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1368 <= _mul_31_source_stop;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1369 <= _tmp_1368;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1370 <= _tmp_1369;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1371 <= _tmp_1370;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1372 <= _tmp_1371;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1373 <= _tmp_1372;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1374 <= _tmp_1373;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1375 <= _tmp_1374;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1376 <= _tmp_1375;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1377 <= _tmp_1376;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1378 <= _mul_31_source_busy;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1379 <= _tmp_1378;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1380 <= _tmp_1379;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1381 <= _tmp_1380;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1382 <= _tmp_1381;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1383 <= _tmp_1382;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1384 <= _tmp_1383;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1385 <= _tmp_1384;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1386 <= _tmp_1385;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1387 <= _tmp_1386;
      end 
      if(_mul_31_stream_oready) begin
        _tmp_1388 <= _mul_31_sink_busy;
      end 
      if(!_mul_31_sink_busy && _tmp_1388) begin
        _mul_31_busy_reg <= 0;
      end 
      if(_mul_31_source_busy) begin
        _mul_31_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_31_fsm_1 = 1;
  localparam _mul_31_fsm_2 = 2;
  localparam _mul_31_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_31_fsm <= _mul_31_fsm_init;
      _mul_31_source_start <= 0;
      _mul_31_source_busy <= 0;
      _mul_31_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_31_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_31_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_31_stream_oready && _tmp_1357) begin
        _mul_31_stream_ivalid <= 1;
      end 
      if(_mul_31_stream_oready && 1'd0) begin
        _mul_31_stream_ivalid <= 0;
      end 
      case(_mul_31_fsm)
        _mul_31_fsm_init: begin
          if(_mul_31_run_flag) begin
            _mul_31_source_start <= 1;
          end 
          if(_mul_31_run_flag) begin
            _mul_31_fsm <= _mul_31_fsm_1;
          end 
        end
        _mul_31_fsm_1: begin
          if(_mul_31_source_start && _mul_31_stream_oready) begin
            _mul_31_source_start <= 0;
            _mul_31_source_busy <= 1;
          end 
          if(_mul_31_source_start && _mul_31_stream_oready) begin
            _mul_31_fsm <= _mul_31_fsm_2;
          end 
        end
        _mul_31_fsm_2: begin
          if(_mul_31_stream_oready) begin
            _mul_31_fsm <= _mul_31_fsm_3;
          end 
        end
        _mul_31_fsm_3: begin
          if(_mul_31_stream_oready && 1'd0) begin
            _mul_31_source_busy <= 0;
          end 
          if(_mul_31_stream_oready && 1'd0 && _mul_31_run_flag) begin
            _mul_31_source_start <= 1;
          end 
          if(_mul_31_stream_oready && 1'd0) begin
            _mul_31_fsm <= _mul_31_fsm_init;
          end 
          if(_mul_31_stream_oready && 1'd0 && _mul_31_run_flag) begin
            _mul_31_fsm <= _mul_31_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_32_x_source_ram_renable <= 0;
      _mul_32_x_source_fifo_deq <= 0;
      _mul_32_x_idle <= 1;
      _mul_32_y_source_ram_renable <= 0;
      _mul_32_y_source_fifo_deq <= 0;
      _mul_32_y_idle <= 1;
      _mul_32_rshift_source_ram_renable <= 0;
      _mul_32_rshift_source_fifo_deq <= 0;
      _mul_32_rshift_idle <= 1;
      _mul_32_z_sink_wenable <= 0;
      _mul_32_z_sink_fifo_enq <= 0;
      __mul_32_stream_ivalid_1 <= 0;
      __mul_32_stream_ivalid_2 <= 0;
      __mul_32_stream_ivalid_3 <= 0;
      __mul_32_stream_ivalid_4 <= 0;
      __mul_32_stream_ivalid_5 <= 0;
      __mul_32_stream_ivalid_6 <= 0;
      __mul_32_stream_ivalid_7 <= 0;
      __mul_32_stream_ivalid_8 <= 0;
      _greaterthan_data_683 <= 0;
      _minus_data_685 <= 0;
      _greatereq_data_696 <= 0;
      __delay_data_2134__variable_680 <= 0;
      __delay_data_2137__variable_681 <= 0;
      __delay_data_2140__variable_682 <= 0;
      _sll_data_687 <= 0;
      __delay_data_2131_greaterthan_683 <= 0;
      __delay_data_2132_greatereq_696 <= 0;
      __delay_data_2135__delay_2134__variable_680 <= 0;
      __delay_data_2138__delay_2137__variable_681 <= 0;
      __delay_data_2141__delay_2140__variable_682 <= 0;
      _cond_data_693 <= 0;
      __delay_data_2133__delay_2132_greatereq_696 <= 0;
      __delay_data_2136__delay_2135__delay_2134__variable_680 <= 0;
      __delay_data_2139__delay_2138__delay_2137__variable_681 <= 0;
      __delay_data_2142__delay_2141__delay_2140__variable_682 <= 0;
      __muladd_madd_odata_reg_699 <= 0;
      __delay_data_2143__delay_2142__delay_2141____variable_682 <= 0;
      __delay_data_2144__delay_2143__delay_2142____variable_682 <= 0;
      __delay_data_2145__delay_2144__delay_2143____variable_682 <= 0;
      __delay_data_2146__delay_2145__delay_2144____variable_682 <= 0;
      _sra_data_700 <= 0;
      __variable_wdata_680 <= 0;
      __variable_wdata_681 <= 0;
      __variable_wdata_682 <= 0;
      _tmp_1389 <= 0;
      _tmp_1390 <= 0;
      _tmp_1391 <= 0;
      _tmp_1392 <= 0;
      _tmp_1393 <= 0;
      _tmp_1394 <= 0;
      _tmp_1395 <= 0;
      _tmp_1396 <= 0;
      _tmp_1397 <= 0;
      _tmp_1398 <= 0;
      _tmp_1399 <= 0;
      _tmp_1400 <= 0;
      _tmp_1401 <= 0;
      _tmp_1402 <= 0;
      _tmp_1403 <= 0;
      _tmp_1404 <= 0;
      _tmp_1405 <= 0;
      _tmp_1406 <= 0;
      _tmp_1407 <= 0;
      _tmp_1408 <= 0;
      _tmp_1409 <= 0;
      _tmp_1410 <= 0;
      _tmp_1411 <= 0;
      _tmp_1412 <= 0;
      _tmp_1413 <= 0;
      _tmp_1414 <= 0;
      _tmp_1415 <= 0;
      _tmp_1416 <= 0;
      _tmp_1417 <= 0;
      _tmp_1418 <= 0;
      _tmp_1419 <= 0;
      _tmp_1420 <= 0;
      _tmp_1421 <= 0;
      _tmp_1422 <= 0;
      _mul_32_busy_reg <= 0;
    end else begin
      if(_mul_32_stream_oready) begin
        _mul_32_x_source_ram_renable <= 0;
        _mul_32_x_source_fifo_deq <= 0;
      end 
      _mul_32_x_idle <= _mul_32_x_idle;
      if(_mul_32_stream_oready) begin
        _mul_32_y_source_ram_renable <= 0;
        _mul_32_y_source_fifo_deq <= 0;
      end 
      _mul_32_y_idle <= _mul_32_y_idle;
      if(_mul_32_stream_oready) begin
        _mul_32_rshift_source_ram_renable <= 0;
        _mul_32_rshift_source_fifo_deq <= 0;
      end 
      _mul_32_rshift_idle <= _mul_32_rshift_idle;
      if(_mul_32_stream_oready) begin
        _mul_32_z_sink_wenable <= 0;
        _mul_32_z_sink_fifo_enq <= 0;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_1 <= _mul_32_stream_ivalid;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_2 <= __mul_32_stream_ivalid_1;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_3 <= __mul_32_stream_ivalid_2;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_4 <= __mul_32_stream_ivalid_3;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_5 <= __mul_32_stream_ivalid_4;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_6 <= __mul_32_stream_ivalid_5;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_7 <= __mul_32_stream_ivalid_6;
      end 
      if(_mul_32_stream_oready) begin
        __mul_32_stream_ivalid_8 <= __mul_32_stream_ivalid_7;
      end 
      if(_mul_32_stream_oready) begin
        _greaterthan_data_683 <= mul_32_rshift_data > 1'sd0;
      end 
      if(_mul_32_stream_oready) begin
        _minus_data_685 <= mul_32_rshift_data - 2'sd1;
      end 
      if(_mul_32_stream_oready) begin
        _greatereq_data_696 <= mul_32_x_data >= 1'sd0;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2134__variable_680 <= mul_32_x_data;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2137__variable_681 <= mul_32_y_data;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2140__variable_682 <= mul_32_rshift_data;
      end 
      if(_mul_32_stream_oready) begin
        _sll_data_687 <= 2'sd1 << _minus_data_685;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2131_greaterthan_683 <= _greaterthan_data_683;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2132_greatereq_696 <= _greatereq_data_696;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2135__delay_2134__variable_680 <= __delay_data_2134__variable_680;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2138__delay_2137__variable_681 <= __delay_data_2137__variable_681;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2141__delay_2140__variable_682 <= __delay_data_2140__variable_682;
      end 
      if(_mul_32_stream_oready) begin
        _cond_data_693 <= (__delay_data_2131_greaterthan_683)? _sll_data_687 : 1'sd0;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2133__delay_2132_greatereq_696 <= __delay_data_2132_greatereq_696;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2136__delay_2135__delay_2134__variable_680 <= __delay_data_2135__delay_2134__variable_680;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2139__delay_2138__delay_2137__variable_681 <= __delay_data_2138__delay_2137__variable_681;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2142__delay_2141__delay_2140__variable_682 <= __delay_data_2141__delay_2140__variable_682;
      end 
      if(_mul_32_stream_oready) begin
        __muladd_madd_odata_reg_699 <= __muladd_madd_odata_699;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2143__delay_2142__delay_2141____variable_682 <= __delay_data_2142__delay_2141__delay_2140__variable_682;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2144__delay_2143__delay_2142____variable_682 <= __delay_data_2143__delay_2142__delay_2141____variable_682;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2145__delay_2144__delay_2143____variable_682 <= __delay_data_2144__delay_2143__delay_2142____variable_682;
      end 
      if(_mul_32_stream_oready) begin
        __delay_data_2146__delay_2145__delay_2144____variable_682 <= __delay_data_2145__delay_2144__delay_2143____variable_682;
      end 
      if(_mul_32_stream_oready) begin
        _sra_data_700 <= __muladd_data_699 >>> __delay_data_2146__delay_2145__delay_2144____variable_682;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_680 <= _cond_data_2011;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_681 <= _cond_data_1539;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_682 <= __delay_data_2919__delay_2918_plus_2147;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1389 <= _mul_32_source_start;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1390 <= _tmp_1389;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1391 <= _tmp_1390;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1392 <= _mul_32_source_start;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1393 <= _tmp_1392;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1394 <= _tmp_1393;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1395 <= _tmp_1394;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1396 <= _tmp_1395;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1397 <= _tmp_1396;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1398 <= _tmp_1397;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1399 <= _tmp_1398;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1400 <= _tmp_1399;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1401 <= _tmp_1400;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1402 <= _mul_32_source_stop;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1403 <= _tmp_1402;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1404 <= _tmp_1403;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1405 <= _tmp_1404;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1406 <= _tmp_1405;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1407 <= _tmp_1406;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1408 <= _tmp_1407;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1409 <= _tmp_1408;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1410 <= _tmp_1409;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1411 <= _tmp_1410;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1412 <= _mul_32_source_busy;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1413 <= _tmp_1412;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1414 <= _tmp_1413;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1415 <= _tmp_1414;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1416 <= _tmp_1415;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1417 <= _tmp_1416;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1418 <= _tmp_1417;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1419 <= _tmp_1418;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1420 <= _tmp_1419;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1421 <= _tmp_1420;
      end 
      if(_mul_32_stream_oready) begin
        _tmp_1422 <= _mul_32_sink_busy;
      end 
      if(!_mul_32_sink_busy && _tmp_1422) begin
        _mul_32_busy_reg <= 0;
      end 
      if(_mul_32_source_busy) begin
        _mul_32_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_32_fsm_1 = 1;
  localparam _mul_32_fsm_2 = 2;
  localparam _mul_32_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_32_fsm <= _mul_32_fsm_init;
      _mul_32_source_start <= 0;
      _mul_32_source_busy <= 0;
      _mul_32_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_32_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_32_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_32_stream_oready && _tmp_1391) begin
        _mul_32_stream_ivalid <= 1;
      end 
      if(_mul_32_stream_oready && 1'd0) begin
        _mul_32_stream_ivalid <= 0;
      end 
      case(_mul_32_fsm)
        _mul_32_fsm_init: begin
          if(_mul_32_run_flag) begin
            _mul_32_source_start <= 1;
          end 
          if(_mul_32_run_flag) begin
            _mul_32_fsm <= _mul_32_fsm_1;
          end 
        end
        _mul_32_fsm_1: begin
          if(_mul_32_source_start && _mul_32_stream_oready) begin
            _mul_32_source_start <= 0;
            _mul_32_source_busy <= 1;
          end 
          if(_mul_32_source_start && _mul_32_stream_oready) begin
            _mul_32_fsm <= _mul_32_fsm_2;
          end 
        end
        _mul_32_fsm_2: begin
          if(_mul_32_stream_oready) begin
            _mul_32_fsm <= _mul_32_fsm_3;
          end 
        end
        _mul_32_fsm_3: begin
          if(_mul_32_stream_oready && 1'd0) begin
            _mul_32_source_busy <= 0;
          end 
          if(_mul_32_stream_oready && 1'd0 && _mul_32_run_flag) begin
            _mul_32_source_start <= 1;
          end 
          if(_mul_32_stream_oready && 1'd0) begin
            _mul_32_fsm <= _mul_32_fsm_init;
          end 
          if(_mul_32_stream_oready && 1'd0 && _mul_32_run_flag) begin
            _mul_32_fsm <= _mul_32_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_33_x_source_ram_renable <= 0;
      _mul_33_x_source_fifo_deq <= 0;
      _mul_33_x_idle <= 1;
      _mul_33_y_source_ram_renable <= 0;
      _mul_33_y_source_fifo_deq <= 0;
      _mul_33_y_idle <= 1;
      _mul_33_rshift_source_ram_renable <= 0;
      _mul_33_rshift_source_fifo_deq <= 0;
      _mul_33_rshift_idle <= 1;
      _mul_33_z_sink_wenable <= 0;
      _mul_33_z_sink_fifo_enq <= 0;
      __mul_33_stream_ivalid_1 <= 0;
      __mul_33_stream_ivalid_2 <= 0;
      __mul_33_stream_ivalid_3 <= 0;
      __mul_33_stream_ivalid_4 <= 0;
      __mul_33_stream_ivalid_5 <= 0;
      __mul_33_stream_ivalid_6 <= 0;
      __mul_33_stream_ivalid_7 <= 0;
      __mul_33_stream_ivalid_8 <= 0;
      _greaterthan_data_704 <= 0;
      _minus_data_706 <= 0;
      _greatereq_data_717 <= 0;
      __delay_data_2153__variable_701 <= 0;
      __delay_data_2156__variable_702 <= 0;
      __delay_data_2159__variable_703 <= 0;
      _sll_data_708 <= 0;
      __delay_data_2150_greaterthan_704 <= 0;
      __delay_data_2151_greatereq_717 <= 0;
      __delay_data_2154__delay_2153__variable_701 <= 0;
      __delay_data_2157__delay_2156__variable_702 <= 0;
      __delay_data_2160__delay_2159__variable_703 <= 0;
      _cond_data_714 <= 0;
      __delay_data_2152__delay_2151_greatereq_717 <= 0;
      __delay_data_2155__delay_2154__delay_2153__variable_701 <= 0;
      __delay_data_2158__delay_2157__delay_2156__variable_702 <= 0;
      __delay_data_2161__delay_2160__delay_2159__variable_703 <= 0;
      __muladd_madd_odata_reg_720 <= 0;
      __delay_data_2162__delay_2161__delay_2160____variable_703 <= 0;
      __delay_data_2163__delay_2162__delay_2161____variable_703 <= 0;
      __delay_data_2164__delay_2163__delay_2162____variable_703 <= 0;
      __delay_data_2165__delay_2164__delay_2163____variable_703 <= 0;
      _sra_data_721 <= 0;
      __variable_wdata_701 <= 0;
      __variable_wdata_702 <= 0;
      __variable_wdata_703 <= 0;
      _tmp_1423 <= 0;
      _tmp_1424 <= 0;
      _tmp_1425 <= 0;
      _tmp_1426 <= 0;
      _tmp_1427 <= 0;
      _tmp_1428 <= 0;
      _tmp_1429 <= 0;
      _tmp_1430 <= 0;
      _tmp_1431 <= 0;
      _tmp_1432 <= 0;
      _tmp_1433 <= 0;
      _tmp_1434 <= 0;
      _tmp_1435 <= 0;
      _tmp_1436 <= 0;
      _tmp_1437 <= 0;
      _tmp_1438 <= 0;
      _tmp_1439 <= 0;
      _tmp_1440 <= 0;
      _tmp_1441 <= 0;
      _tmp_1442 <= 0;
      _tmp_1443 <= 0;
      _tmp_1444 <= 0;
      _tmp_1445 <= 0;
      _tmp_1446 <= 0;
      _tmp_1447 <= 0;
      _tmp_1448 <= 0;
      _tmp_1449 <= 0;
      _tmp_1450 <= 0;
      _tmp_1451 <= 0;
      _tmp_1452 <= 0;
      _tmp_1453 <= 0;
      _tmp_1454 <= 0;
      _tmp_1455 <= 0;
      _tmp_1456 <= 0;
      _mul_33_busy_reg <= 0;
    end else begin
      if(_mul_33_stream_oready) begin
        _mul_33_x_source_ram_renable <= 0;
        _mul_33_x_source_fifo_deq <= 0;
      end 
      _mul_33_x_idle <= _mul_33_x_idle;
      if(_mul_33_stream_oready) begin
        _mul_33_y_source_ram_renable <= 0;
        _mul_33_y_source_fifo_deq <= 0;
      end 
      _mul_33_y_idle <= _mul_33_y_idle;
      if(_mul_33_stream_oready) begin
        _mul_33_rshift_source_ram_renable <= 0;
        _mul_33_rshift_source_fifo_deq <= 0;
      end 
      _mul_33_rshift_idle <= _mul_33_rshift_idle;
      if(_mul_33_stream_oready) begin
        _mul_33_z_sink_wenable <= 0;
        _mul_33_z_sink_fifo_enq <= 0;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_1 <= _mul_33_stream_ivalid;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_2 <= __mul_33_stream_ivalid_1;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_3 <= __mul_33_stream_ivalid_2;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_4 <= __mul_33_stream_ivalid_3;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_5 <= __mul_33_stream_ivalid_4;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_6 <= __mul_33_stream_ivalid_5;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_7 <= __mul_33_stream_ivalid_6;
      end 
      if(_mul_33_stream_oready) begin
        __mul_33_stream_ivalid_8 <= __mul_33_stream_ivalid_7;
      end 
      if(_mul_33_stream_oready) begin
        _greaterthan_data_704 <= mul_33_rshift_data > 1'sd0;
      end 
      if(_mul_33_stream_oready) begin
        _minus_data_706 <= mul_33_rshift_data - 2'sd1;
      end 
      if(_mul_33_stream_oready) begin
        _greatereq_data_717 <= mul_33_x_data >= 1'sd0;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2153__variable_701 <= mul_33_x_data;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2156__variable_702 <= mul_33_y_data;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2159__variable_703 <= mul_33_rshift_data;
      end 
      if(_mul_33_stream_oready) begin
        _sll_data_708 <= 2'sd1 << _minus_data_706;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2150_greaterthan_704 <= _greaterthan_data_704;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2151_greatereq_717 <= _greatereq_data_717;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2154__delay_2153__variable_701 <= __delay_data_2153__variable_701;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2157__delay_2156__variable_702 <= __delay_data_2156__variable_702;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2160__delay_2159__variable_703 <= __delay_data_2159__variable_703;
      end 
      if(_mul_33_stream_oready) begin
        _cond_data_714 <= (__delay_data_2150_greaterthan_704)? _sll_data_708 : 1'sd0;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2152__delay_2151_greatereq_717 <= __delay_data_2151_greatereq_717;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2155__delay_2154__delay_2153__variable_701 <= __delay_data_2154__delay_2153__variable_701;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2158__delay_2157__delay_2156__variable_702 <= __delay_data_2157__delay_2156__variable_702;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2161__delay_2160__delay_2159__variable_703 <= __delay_data_2160__delay_2159__variable_703;
      end 
      if(_mul_33_stream_oready) begin
        __muladd_madd_odata_reg_720 <= __muladd_madd_odata_720;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2162__delay_2161__delay_2160____variable_703 <= __delay_data_2161__delay_2160__delay_2159__variable_703;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2163__delay_2162__delay_2161____variable_703 <= __delay_data_2162__delay_2161__delay_2160____variable_703;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2164__delay_2163__delay_2162____variable_703 <= __delay_data_2163__delay_2162__delay_2161____variable_703;
      end 
      if(_mul_33_stream_oready) begin
        __delay_data_2165__delay_2164__delay_2163____variable_703 <= __delay_data_2164__delay_2163__delay_2162____variable_703;
      end 
      if(_mul_33_stream_oready) begin
        _sra_data_721 <= __muladd_data_720 >>> __delay_data_2165__delay_2164__delay_2163____variable_703;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_701 <= _cond_data_2013;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_702 <= _cond_data_1541;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_703 <= __delay_data_2929__delay_2928_plus_2166;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1423 <= _mul_33_source_start;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1424 <= _tmp_1423;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1425 <= _tmp_1424;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1426 <= _mul_33_source_start;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1427 <= _tmp_1426;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1428 <= _tmp_1427;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1429 <= _tmp_1428;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1430 <= _tmp_1429;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1431 <= _tmp_1430;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1432 <= _tmp_1431;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1433 <= _tmp_1432;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1434 <= _tmp_1433;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1435 <= _tmp_1434;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1436 <= _mul_33_source_stop;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1437 <= _tmp_1436;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1438 <= _tmp_1437;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1439 <= _tmp_1438;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1440 <= _tmp_1439;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1441 <= _tmp_1440;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1442 <= _tmp_1441;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1443 <= _tmp_1442;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1444 <= _tmp_1443;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1445 <= _tmp_1444;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1446 <= _mul_33_source_busy;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1447 <= _tmp_1446;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1448 <= _tmp_1447;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1449 <= _tmp_1448;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1450 <= _tmp_1449;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1451 <= _tmp_1450;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1452 <= _tmp_1451;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1453 <= _tmp_1452;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1454 <= _tmp_1453;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1455 <= _tmp_1454;
      end 
      if(_mul_33_stream_oready) begin
        _tmp_1456 <= _mul_33_sink_busy;
      end 
      if(!_mul_33_sink_busy && _tmp_1456) begin
        _mul_33_busy_reg <= 0;
      end 
      if(_mul_33_source_busy) begin
        _mul_33_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_33_fsm_1 = 1;
  localparam _mul_33_fsm_2 = 2;
  localparam _mul_33_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_33_fsm <= _mul_33_fsm_init;
      _mul_33_source_start <= 0;
      _mul_33_source_busy <= 0;
      _mul_33_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_33_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_33_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_33_stream_oready && _tmp_1425) begin
        _mul_33_stream_ivalid <= 1;
      end 
      if(_mul_33_stream_oready && 1'd0) begin
        _mul_33_stream_ivalid <= 0;
      end 
      case(_mul_33_fsm)
        _mul_33_fsm_init: begin
          if(_mul_33_run_flag) begin
            _mul_33_source_start <= 1;
          end 
          if(_mul_33_run_flag) begin
            _mul_33_fsm <= _mul_33_fsm_1;
          end 
        end
        _mul_33_fsm_1: begin
          if(_mul_33_source_start && _mul_33_stream_oready) begin
            _mul_33_source_start <= 0;
            _mul_33_source_busy <= 1;
          end 
          if(_mul_33_source_start && _mul_33_stream_oready) begin
            _mul_33_fsm <= _mul_33_fsm_2;
          end 
        end
        _mul_33_fsm_2: begin
          if(_mul_33_stream_oready) begin
            _mul_33_fsm <= _mul_33_fsm_3;
          end 
        end
        _mul_33_fsm_3: begin
          if(_mul_33_stream_oready && 1'd0) begin
            _mul_33_source_busy <= 0;
          end 
          if(_mul_33_stream_oready && 1'd0 && _mul_33_run_flag) begin
            _mul_33_source_start <= 1;
          end 
          if(_mul_33_stream_oready && 1'd0) begin
            _mul_33_fsm <= _mul_33_fsm_init;
          end 
          if(_mul_33_stream_oready && 1'd0 && _mul_33_run_flag) begin
            _mul_33_fsm <= _mul_33_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_34_x_source_ram_renable <= 0;
      _mul_34_x_source_fifo_deq <= 0;
      _mul_34_x_idle <= 1;
      _mul_34_y_source_ram_renable <= 0;
      _mul_34_y_source_fifo_deq <= 0;
      _mul_34_y_idle <= 1;
      _mul_34_rshift_source_ram_renable <= 0;
      _mul_34_rshift_source_fifo_deq <= 0;
      _mul_34_rshift_idle <= 1;
      _mul_34_z_sink_wenable <= 0;
      _mul_34_z_sink_fifo_enq <= 0;
      __mul_34_stream_ivalid_1 <= 0;
      __mul_34_stream_ivalid_2 <= 0;
      __mul_34_stream_ivalid_3 <= 0;
      __mul_34_stream_ivalid_4 <= 0;
      __mul_34_stream_ivalid_5 <= 0;
      __mul_34_stream_ivalid_6 <= 0;
      __mul_34_stream_ivalid_7 <= 0;
      __mul_34_stream_ivalid_8 <= 0;
      _greaterthan_data_725 <= 0;
      _minus_data_727 <= 0;
      _greatereq_data_738 <= 0;
      __delay_data_2172__variable_722 <= 0;
      __delay_data_2175__variable_723 <= 0;
      __delay_data_2178__variable_724 <= 0;
      _sll_data_729 <= 0;
      __delay_data_2169_greaterthan_725 <= 0;
      __delay_data_2170_greatereq_738 <= 0;
      __delay_data_2173__delay_2172__variable_722 <= 0;
      __delay_data_2176__delay_2175__variable_723 <= 0;
      __delay_data_2179__delay_2178__variable_724 <= 0;
      _cond_data_735 <= 0;
      __delay_data_2171__delay_2170_greatereq_738 <= 0;
      __delay_data_2174__delay_2173__delay_2172__variable_722 <= 0;
      __delay_data_2177__delay_2176__delay_2175__variable_723 <= 0;
      __delay_data_2180__delay_2179__delay_2178__variable_724 <= 0;
      __muladd_madd_odata_reg_741 <= 0;
      __delay_data_2181__delay_2180__delay_2179____variable_724 <= 0;
      __delay_data_2182__delay_2181__delay_2180____variable_724 <= 0;
      __delay_data_2183__delay_2182__delay_2181____variable_724 <= 0;
      __delay_data_2184__delay_2183__delay_2182____variable_724 <= 0;
      _sra_data_742 <= 0;
      __variable_wdata_722 <= 0;
      __variable_wdata_723 <= 0;
      __variable_wdata_724 <= 0;
      _tmp_1457 <= 0;
      _tmp_1458 <= 0;
      _tmp_1459 <= 0;
      _tmp_1460 <= 0;
      _tmp_1461 <= 0;
      _tmp_1462 <= 0;
      _tmp_1463 <= 0;
      _tmp_1464 <= 0;
      _tmp_1465 <= 0;
      _tmp_1466 <= 0;
      _tmp_1467 <= 0;
      _tmp_1468 <= 0;
      _tmp_1469 <= 0;
      _tmp_1470 <= 0;
      _tmp_1471 <= 0;
      _tmp_1472 <= 0;
      _tmp_1473 <= 0;
      _tmp_1474 <= 0;
      _tmp_1475 <= 0;
      _tmp_1476 <= 0;
      _tmp_1477 <= 0;
      _tmp_1478 <= 0;
      _tmp_1479 <= 0;
      _tmp_1480 <= 0;
      _tmp_1481 <= 0;
      _tmp_1482 <= 0;
      _tmp_1483 <= 0;
      _tmp_1484 <= 0;
      _tmp_1485 <= 0;
      _tmp_1486 <= 0;
      _tmp_1487 <= 0;
      _tmp_1488 <= 0;
      _tmp_1489 <= 0;
      _tmp_1490 <= 0;
      _mul_34_busy_reg <= 0;
    end else begin
      if(_mul_34_stream_oready) begin
        _mul_34_x_source_ram_renable <= 0;
        _mul_34_x_source_fifo_deq <= 0;
      end 
      _mul_34_x_idle <= _mul_34_x_idle;
      if(_mul_34_stream_oready) begin
        _mul_34_y_source_ram_renable <= 0;
        _mul_34_y_source_fifo_deq <= 0;
      end 
      _mul_34_y_idle <= _mul_34_y_idle;
      if(_mul_34_stream_oready) begin
        _mul_34_rshift_source_ram_renable <= 0;
        _mul_34_rshift_source_fifo_deq <= 0;
      end 
      _mul_34_rshift_idle <= _mul_34_rshift_idle;
      if(_mul_34_stream_oready) begin
        _mul_34_z_sink_wenable <= 0;
        _mul_34_z_sink_fifo_enq <= 0;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_1 <= _mul_34_stream_ivalid;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_2 <= __mul_34_stream_ivalid_1;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_3 <= __mul_34_stream_ivalid_2;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_4 <= __mul_34_stream_ivalid_3;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_5 <= __mul_34_stream_ivalid_4;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_6 <= __mul_34_stream_ivalid_5;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_7 <= __mul_34_stream_ivalid_6;
      end 
      if(_mul_34_stream_oready) begin
        __mul_34_stream_ivalid_8 <= __mul_34_stream_ivalid_7;
      end 
      if(_mul_34_stream_oready) begin
        _greaterthan_data_725 <= mul_34_rshift_data > 1'sd0;
      end 
      if(_mul_34_stream_oready) begin
        _minus_data_727 <= mul_34_rshift_data - 2'sd1;
      end 
      if(_mul_34_stream_oready) begin
        _greatereq_data_738 <= mul_34_x_data >= 1'sd0;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2172__variable_722 <= mul_34_x_data;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2175__variable_723 <= mul_34_y_data;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2178__variable_724 <= mul_34_rshift_data;
      end 
      if(_mul_34_stream_oready) begin
        _sll_data_729 <= 2'sd1 << _minus_data_727;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2169_greaterthan_725 <= _greaterthan_data_725;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2170_greatereq_738 <= _greatereq_data_738;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2173__delay_2172__variable_722 <= __delay_data_2172__variable_722;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2176__delay_2175__variable_723 <= __delay_data_2175__variable_723;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2179__delay_2178__variable_724 <= __delay_data_2178__variable_724;
      end 
      if(_mul_34_stream_oready) begin
        _cond_data_735 <= (__delay_data_2169_greaterthan_725)? _sll_data_729 : 1'sd0;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2171__delay_2170_greatereq_738 <= __delay_data_2170_greatereq_738;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2174__delay_2173__delay_2172__variable_722 <= __delay_data_2173__delay_2172__variable_722;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2177__delay_2176__delay_2175__variable_723 <= __delay_data_2176__delay_2175__variable_723;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2180__delay_2179__delay_2178__variable_724 <= __delay_data_2179__delay_2178__variable_724;
      end 
      if(_mul_34_stream_oready) begin
        __muladd_madd_odata_reg_741 <= __muladd_madd_odata_741;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2181__delay_2180__delay_2179____variable_724 <= __delay_data_2180__delay_2179__delay_2178__variable_724;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2182__delay_2181__delay_2180____variable_724 <= __delay_data_2181__delay_2180__delay_2179____variable_724;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2183__delay_2182__delay_2181____variable_724 <= __delay_data_2182__delay_2181__delay_2180____variable_724;
      end 
      if(_mul_34_stream_oready) begin
        __delay_data_2184__delay_2183__delay_2182____variable_724 <= __delay_data_2183__delay_2182__delay_2181____variable_724;
      end 
      if(_mul_34_stream_oready) begin
        _sra_data_742 <= __muladd_data_741 >>> __delay_data_2184__delay_2183__delay_2182____variable_724;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_722 <= _cond_data_2015;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_723 <= _cond_data_1543;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_724 <= __delay_data_2939__delay_2938_plus_2185;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1457 <= _mul_34_source_start;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1458 <= _tmp_1457;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1459 <= _tmp_1458;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1460 <= _mul_34_source_start;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1461 <= _tmp_1460;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1462 <= _tmp_1461;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1463 <= _tmp_1462;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1464 <= _tmp_1463;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1465 <= _tmp_1464;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1466 <= _tmp_1465;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1467 <= _tmp_1466;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1468 <= _tmp_1467;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1469 <= _tmp_1468;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1470 <= _mul_34_source_stop;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1471 <= _tmp_1470;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1472 <= _tmp_1471;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1473 <= _tmp_1472;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1474 <= _tmp_1473;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1475 <= _tmp_1474;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1476 <= _tmp_1475;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1477 <= _tmp_1476;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1478 <= _tmp_1477;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1479 <= _tmp_1478;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1480 <= _mul_34_source_busy;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1481 <= _tmp_1480;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1482 <= _tmp_1481;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1483 <= _tmp_1482;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1484 <= _tmp_1483;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1485 <= _tmp_1484;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1486 <= _tmp_1485;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1487 <= _tmp_1486;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1488 <= _tmp_1487;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1489 <= _tmp_1488;
      end 
      if(_mul_34_stream_oready) begin
        _tmp_1490 <= _mul_34_sink_busy;
      end 
      if(!_mul_34_sink_busy && _tmp_1490) begin
        _mul_34_busy_reg <= 0;
      end 
      if(_mul_34_source_busy) begin
        _mul_34_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_34_fsm_1 = 1;
  localparam _mul_34_fsm_2 = 2;
  localparam _mul_34_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_34_fsm <= _mul_34_fsm_init;
      _mul_34_source_start <= 0;
      _mul_34_source_busy <= 0;
      _mul_34_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_34_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_34_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_34_stream_oready && _tmp_1459) begin
        _mul_34_stream_ivalid <= 1;
      end 
      if(_mul_34_stream_oready && 1'd0) begin
        _mul_34_stream_ivalid <= 0;
      end 
      case(_mul_34_fsm)
        _mul_34_fsm_init: begin
          if(_mul_34_run_flag) begin
            _mul_34_source_start <= 1;
          end 
          if(_mul_34_run_flag) begin
            _mul_34_fsm <= _mul_34_fsm_1;
          end 
        end
        _mul_34_fsm_1: begin
          if(_mul_34_source_start && _mul_34_stream_oready) begin
            _mul_34_source_start <= 0;
            _mul_34_source_busy <= 1;
          end 
          if(_mul_34_source_start && _mul_34_stream_oready) begin
            _mul_34_fsm <= _mul_34_fsm_2;
          end 
        end
        _mul_34_fsm_2: begin
          if(_mul_34_stream_oready) begin
            _mul_34_fsm <= _mul_34_fsm_3;
          end 
        end
        _mul_34_fsm_3: begin
          if(_mul_34_stream_oready && 1'd0) begin
            _mul_34_source_busy <= 0;
          end 
          if(_mul_34_stream_oready && 1'd0 && _mul_34_run_flag) begin
            _mul_34_source_start <= 1;
          end 
          if(_mul_34_stream_oready && 1'd0) begin
            _mul_34_fsm <= _mul_34_fsm_init;
          end 
          if(_mul_34_stream_oready && 1'd0 && _mul_34_run_flag) begin
            _mul_34_fsm <= _mul_34_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_35_x_source_ram_renable <= 0;
      _mul_35_x_source_fifo_deq <= 0;
      _mul_35_x_idle <= 1;
      _mul_35_y_source_ram_renable <= 0;
      _mul_35_y_source_fifo_deq <= 0;
      _mul_35_y_idle <= 1;
      _mul_35_rshift_source_ram_renable <= 0;
      _mul_35_rshift_source_fifo_deq <= 0;
      _mul_35_rshift_idle <= 1;
      _mul_35_z_sink_wenable <= 0;
      _mul_35_z_sink_fifo_enq <= 0;
      __mul_35_stream_ivalid_1 <= 0;
      __mul_35_stream_ivalid_2 <= 0;
      __mul_35_stream_ivalid_3 <= 0;
      __mul_35_stream_ivalid_4 <= 0;
      __mul_35_stream_ivalid_5 <= 0;
      __mul_35_stream_ivalid_6 <= 0;
      __mul_35_stream_ivalid_7 <= 0;
      __mul_35_stream_ivalid_8 <= 0;
      _greaterthan_data_746 <= 0;
      _minus_data_748 <= 0;
      _greatereq_data_759 <= 0;
      __delay_data_2209__variable_743 <= 0;
      __delay_data_2212__variable_744 <= 0;
      __delay_data_2215__variable_745 <= 0;
      _sll_data_750 <= 0;
      __delay_data_2206_greaterthan_746 <= 0;
      __delay_data_2207_greatereq_759 <= 0;
      __delay_data_2210__delay_2209__variable_743 <= 0;
      __delay_data_2213__delay_2212__variable_744 <= 0;
      __delay_data_2216__delay_2215__variable_745 <= 0;
      _cond_data_756 <= 0;
      __delay_data_2208__delay_2207_greatereq_759 <= 0;
      __delay_data_2211__delay_2210__delay_2209__variable_743 <= 0;
      __delay_data_2214__delay_2213__delay_2212__variable_744 <= 0;
      __delay_data_2217__delay_2216__delay_2215__variable_745 <= 0;
      __muladd_madd_odata_reg_762 <= 0;
      __delay_data_2218__delay_2217__delay_2216____variable_745 <= 0;
      __delay_data_2219__delay_2218__delay_2217____variable_745 <= 0;
      __delay_data_2220__delay_2219__delay_2218____variable_745 <= 0;
      __delay_data_2221__delay_2220__delay_2219____variable_745 <= 0;
      _sra_data_763 <= 0;
      __variable_wdata_743 <= 0;
      __variable_wdata_744 <= 0;
      __variable_wdata_745 <= 0;
      _tmp_1491 <= 0;
      _tmp_1492 <= 0;
      _tmp_1493 <= 0;
      _tmp_1494 <= 0;
      _tmp_1495 <= 0;
      _tmp_1496 <= 0;
      _tmp_1497 <= 0;
      _tmp_1498 <= 0;
      _tmp_1499 <= 0;
      _tmp_1500 <= 0;
      _tmp_1501 <= 0;
      _tmp_1502 <= 0;
      _tmp_1503 <= 0;
      _tmp_1504 <= 0;
      _tmp_1505 <= 0;
      _tmp_1506 <= 0;
      _tmp_1507 <= 0;
      _tmp_1508 <= 0;
      _tmp_1509 <= 0;
      _tmp_1510 <= 0;
      _tmp_1511 <= 0;
      _tmp_1512 <= 0;
      _tmp_1513 <= 0;
      _tmp_1514 <= 0;
      _tmp_1515 <= 0;
      _tmp_1516 <= 0;
      _tmp_1517 <= 0;
      _tmp_1518 <= 0;
      _tmp_1519 <= 0;
      _tmp_1520 <= 0;
      _tmp_1521 <= 0;
      _tmp_1522 <= 0;
      _tmp_1523 <= 0;
      _tmp_1524 <= 0;
      _mul_35_busy_reg <= 0;
    end else begin
      if(_mul_35_stream_oready) begin
        _mul_35_x_source_ram_renable <= 0;
        _mul_35_x_source_fifo_deq <= 0;
      end 
      _mul_35_x_idle <= _mul_35_x_idle;
      if(_mul_35_stream_oready) begin
        _mul_35_y_source_ram_renable <= 0;
        _mul_35_y_source_fifo_deq <= 0;
      end 
      _mul_35_y_idle <= _mul_35_y_idle;
      if(_mul_35_stream_oready) begin
        _mul_35_rshift_source_ram_renable <= 0;
        _mul_35_rshift_source_fifo_deq <= 0;
      end 
      _mul_35_rshift_idle <= _mul_35_rshift_idle;
      if(_mul_35_stream_oready) begin
        _mul_35_z_sink_wenable <= 0;
        _mul_35_z_sink_fifo_enq <= 0;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_1 <= _mul_35_stream_ivalid;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_2 <= __mul_35_stream_ivalid_1;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_3 <= __mul_35_stream_ivalid_2;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_4 <= __mul_35_stream_ivalid_3;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_5 <= __mul_35_stream_ivalid_4;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_6 <= __mul_35_stream_ivalid_5;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_7 <= __mul_35_stream_ivalid_6;
      end 
      if(_mul_35_stream_oready) begin
        __mul_35_stream_ivalid_8 <= __mul_35_stream_ivalid_7;
      end 
      if(_mul_35_stream_oready) begin
        _greaterthan_data_746 <= mul_35_rshift_data > 1'sd0;
      end 
      if(_mul_35_stream_oready) begin
        _minus_data_748 <= mul_35_rshift_data - 2'sd1;
      end 
      if(_mul_35_stream_oready) begin
        _greatereq_data_759 <= mul_35_x_data >= 1'sd0;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2209__variable_743 <= mul_35_x_data;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2212__variable_744 <= mul_35_y_data;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2215__variable_745 <= mul_35_rshift_data;
      end 
      if(_mul_35_stream_oready) begin
        _sll_data_750 <= 2'sd1 << _minus_data_748;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2206_greaterthan_746 <= _greaterthan_data_746;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2207_greatereq_759 <= _greatereq_data_759;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2210__delay_2209__variable_743 <= __delay_data_2209__variable_743;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2213__delay_2212__variable_744 <= __delay_data_2212__variable_744;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2216__delay_2215__variable_745 <= __delay_data_2215__variable_745;
      end 
      if(_mul_35_stream_oready) begin
        _cond_data_756 <= (__delay_data_2206_greaterthan_746)? _sll_data_750 : 1'sd0;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2208__delay_2207_greatereq_759 <= __delay_data_2207_greatereq_759;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2211__delay_2210__delay_2209__variable_743 <= __delay_data_2210__delay_2209__variable_743;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2214__delay_2213__delay_2212__variable_744 <= __delay_data_2213__delay_2212__variable_744;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2217__delay_2216__delay_2215__variable_745 <= __delay_data_2216__delay_2215__variable_745;
      end 
      if(_mul_35_stream_oready) begin
        __muladd_madd_odata_reg_762 <= __muladd_madd_odata_762;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2218__delay_2217__delay_2216____variable_745 <= __delay_data_2217__delay_2216__delay_2215__variable_745;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2219__delay_2218__delay_2217____variable_745 <= __delay_data_2218__delay_2217__delay_2216____variable_745;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2220__delay_2219__delay_2218____variable_745 <= __delay_data_2219__delay_2218__delay_2217____variable_745;
      end 
      if(_mul_35_stream_oready) begin
        __delay_data_2221__delay_2220__delay_2219____variable_745 <= __delay_data_2220__delay_2219__delay_2218____variable_745;
      end 
      if(_mul_35_stream_oready) begin
        _sra_data_763 <= __muladd_data_762 >>> __delay_data_2221__delay_2220__delay_2219____variable_745;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_743 <= _cond_data_2188;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_744 <= _cond_data_1545;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_745 <= __delay_data_2864__delay_2863_plus_2222;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1491 <= _mul_35_source_start;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1492 <= _tmp_1491;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1493 <= _tmp_1492;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1494 <= _mul_35_source_start;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1495 <= _tmp_1494;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1496 <= _tmp_1495;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1497 <= _tmp_1496;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1498 <= _tmp_1497;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1499 <= _tmp_1498;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1500 <= _tmp_1499;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1501 <= _tmp_1500;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1502 <= _tmp_1501;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1503 <= _tmp_1502;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1504 <= _mul_35_source_stop;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1505 <= _tmp_1504;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1506 <= _tmp_1505;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1507 <= _tmp_1506;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1508 <= _tmp_1507;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1509 <= _tmp_1508;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1510 <= _tmp_1509;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1511 <= _tmp_1510;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1512 <= _tmp_1511;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1513 <= _tmp_1512;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1514 <= _mul_35_source_busy;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1515 <= _tmp_1514;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1516 <= _tmp_1515;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1517 <= _tmp_1516;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1518 <= _tmp_1517;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1519 <= _tmp_1518;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1520 <= _tmp_1519;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1521 <= _tmp_1520;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1522 <= _tmp_1521;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1523 <= _tmp_1522;
      end 
      if(_mul_35_stream_oready) begin
        _tmp_1524 <= _mul_35_sink_busy;
      end 
      if(!_mul_35_sink_busy && _tmp_1524) begin
        _mul_35_busy_reg <= 0;
      end 
      if(_mul_35_source_busy) begin
        _mul_35_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_35_fsm_1 = 1;
  localparam _mul_35_fsm_2 = 2;
  localparam _mul_35_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_35_fsm <= _mul_35_fsm_init;
      _mul_35_source_start <= 0;
      _mul_35_source_busy <= 0;
      _mul_35_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_35_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_35_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_35_stream_oready && _tmp_1493) begin
        _mul_35_stream_ivalid <= 1;
      end 
      if(_mul_35_stream_oready && 1'd0) begin
        _mul_35_stream_ivalid <= 0;
      end 
      case(_mul_35_fsm)
        _mul_35_fsm_init: begin
          if(_mul_35_run_flag) begin
            _mul_35_source_start <= 1;
          end 
          if(_mul_35_run_flag) begin
            _mul_35_fsm <= _mul_35_fsm_1;
          end 
        end
        _mul_35_fsm_1: begin
          if(_mul_35_source_start && _mul_35_stream_oready) begin
            _mul_35_source_start <= 0;
            _mul_35_source_busy <= 1;
          end 
          if(_mul_35_source_start && _mul_35_stream_oready) begin
            _mul_35_fsm <= _mul_35_fsm_2;
          end 
        end
        _mul_35_fsm_2: begin
          if(_mul_35_stream_oready) begin
            _mul_35_fsm <= _mul_35_fsm_3;
          end 
        end
        _mul_35_fsm_3: begin
          if(_mul_35_stream_oready && 1'd0) begin
            _mul_35_source_busy <= 0;
          end 
          if(_mul_35_stream_oready && 1'd0 && _mul_35_run_flag) begin
            _mul_35_source_start <= 1;
          end 
          if(_mul_35_stream_oready && 1'd0) begin
            _mul_35_fsm <= _mul_35_fsm_init;
          end 
          if(_mul_35_stream_oready && 1'd0 && _mul_35_run_flag) begin
            _mul_35_fsm <= _mul_35_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_36_x_source_ram_renable <= 0;
      _mul_36_x_source_fifo_deq <= 0;
      _mul_36_x_idle <= 1;
      _mul_36_y_source_ram_renable <= 0;
      _mul_36_y_source_fifo_deq <= 0;
      _mul_36_y_idle <= 1;
      _mul_36_rshift_source_ram_renable <= 0;
      _mul_36_rshift_source_fifo_deq <= 0;
      _mul_36_rshift_idle <= 1;
      _mul_36_z_sink_wenable <= 0;
      _mul_36_z_sink_fifo_enq <= 0;
      __mul_36_stream_ivalid_1 <= 0;
      __mul_36_stream_ivalid_2 <= 0;
      __mul_36_stream_ivalid_3 <= 0;
      __mul_36_stream_ivalid_4 <= 0;
      __mul_36_stream_ivalid_5 <= 0;
      __mul_36_stream_ivalid_6 <= 0;
      __mul_36_stream_ivalid_7 <= 0;
      __mul_36_stream_ivalid_8 <= 0;
      _greaterthan_data_767 <= 0;
      _minus_data_769 <= 0;
      _greatereq_data_780 <= 0;
      __delay_data_2228__variable_764 <= 0;
      __delay_data_2231__variable_765 <= 0;
      __delay_data_2234__variable_766 <= 0;
      _sll_data_771 <= 0;
      __delay_data_2225_greaterthan_767 <= 0;
      __delay_data_2226_greatereq_780 <= 0;
      __delay_data_2229__delay_2228__variable_764 <= 0;
      __delay_data_2232__delay_2231__variable_765 <= 0;
      __delay_data_2235__delay_2234__variable_766 <= 0;
      _cond_data_777 <= 0;
      __delay_data_2227__delay_2226_greatereq_780 <= 0;
      __delay_data_2230__delay_2229__delay_2228__variable_764 <= 0;
      __delay_data_2233__delay_2232__delay_2231__variable_765 <= 0;
      __delay_data_2236__delay_2235__delay_2234__variable_766 <= 0;
      __muladd_madd_odata_reg_783 <= 0;
      __delay_data_2237__delay_2236__delay_2235____variable_766 <= 0;
      __delay_data_2238__delay_2237__delay_2236____variable_766 <= 0;
      __delay_data_2239__delay_2238__delay_2237____variable_766 <= 0;
      __delay_data_2240__delay_2239__delay_2238____variable_766 <= 0;
      _sra_data_784 <= 0;
      __variable_wdata_764 <= 0;
      __variable_wdata_765 <= 0;
      __variable_wdata_766 <= 0;
      _tmp_1525 <= 0;
      _tmp_1526 <= 0;
      _tmp_1527 <= 0;
      _tmp_1528 <= 0;
      _tmp_1529 <= 0;
      _tmp_1530 <= 0;
      _tmp_1531 <= 0;
      _tmp_1532 <= 0;
      _tmp_1533 <= 0;
      _tmp_1534 <= 0;
      _tmp_1535 <= 0;
      _tmp_1536 <= 0;
      _tmp_1537 <= 0;
      _tmp_1538 <= 0;
      _tmp_1539 <= 0;
      _tmp_1540 <= 0;
      _tmp_1541 <= 0;
      _tmp_1542 <= 0;
      _tmp_1543 <= 0;
      _tmp_1544 <= 0;
      _tmp_1545 <= 0;
      _tmp_1546 <= 0;
      _tmp_1547 <= 0;
      _tmp_1548 <= 0;
      _tmp_1549 <= 0;
      _tmp_1550 <= 0;
      _tmp_1551 <= 0;
      _tmp_1552 <= 0;
      _tmp_1553 <= 0;
      _tmp_1554 <= 0;
      _tmp_1555 <= 0;
      _tmp_1556 <= 0;
      _tmp_1557 <= 0;
      _tmp_1558 <= 0;
      _mul_36_busy_reg <= 0;
    end else begin
      if(_mul_36_stream_oready) begin
        _mul_36_x_source_ram_renable <= 0;
        _mul_36_x_source_fifo_deq <= 0;
      end 
      _mul_36_x_idle <= _mul_36_x_idle;
      if(_mul_36_stream_oready) begin
        _mul_36_y_source_ram_renable <= 0;
        _mul_36_y_source_fifo_deq <= 0;
      end 
      _mul_36_y_idle <= _mul_36_y_idle;
      if(_mul_36_stream_oready) begin
        _mul_36_rshift_source_ram_renable <= 0;
        _mul_36_rshift_source_fifo_deq <= 0;
      end 
      _mul_36_rshift_idle <= _mul_36_rshift_idle;
      if(_mul_36_stream_oready) begin
        _mul_36_z_sink_wenable <= 0;
        _mul_36_z_sink_fifo_enq <= 0;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_1 <= _mul_36_stream_ivalid;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_2 <= __mul_36_stream_ivalid_1;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_3 <= __mul_36_stream_ivalid_2;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_4 <= __mul_36_stream_ivalid_3;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_5 <= __mul_36_stream_ivalid_4;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_6 <= __mul_36_stream_ivalid_5;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_7 <= __mul_36_stream_ivalid_6;
      end 
      if(_mul_36_stream_oready) begin
        __mul_36_stream_ivalid_8 <= __mul_36_stream_ivalid_7;
      end 
      if(_mul_36_stream_oready) begin
        _greaterthan_data_767 <= mul_36_rshift_data > 1'sd0;
      end 
      if(_mul_36_stream_oready) begin
        _minus_data_769 <= mul_36_rshift_data - 2'sd1;
      end 
      if(_mul_36_stream_oready) begin
        _greatereq_data_780 <= mul_36_x_data >= 1'sd0;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2228__variable_764 <= mul_36_x_data;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2231__variable_765 <= mul_36_y_data;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2234__variable_766 <= mul_36_rshift_data;
      end 
      if(_mul_36_stream_oready) begin
        _sll_data_771 <= 2'sd1 << _minus_data_769;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2225_greaterthan_767 <= _greaterthan_data_767;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2226_greatereq_780 <= _greatereq_data_780;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2229__delay_2228__variable_764 <= __delay_data_2228__variable_764;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2232__delay_2231__variable_765 <= __delay_data_2231__variable_765;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2235__delay_2234__variable_766 <= __delay_data_2234__variable_766;
      end 
      if(_mul_36_stream_oready) begin
        _cond_data_777 <= (__delay_data_2225_greaterthan_767)? _sll_data_771 : 1'sd0;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2227__delay_2226_greatereq_780 <= __delay_data_2226_greatereq_780;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2230__delay_2229__delay_2228__variable_764 <= __delay_data_2229__delay_2228__variable_764;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2233__delay_2232__delay_2231__variable_765 <= __delay_data_2232__delay_2231__variable_765;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2236__delay_2235__delay_2234__variable_766 <= __delay_data_2235__delay_2234__variable_766;
      end 
      if(_mul_36_stream_oready) begin
        __muladd_madd_odata_reg_783 <= __muladd_madd_odata_783;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2237__delay_2236__delay_2235____variable_766 <= __delay_data_2236__delay_2235__delay_2234__variable_766;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2238__delay_2237__delay_2236____variable_766 <= __delay_data_2237__delay_2236__delay_2235____variable_766;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2239__delay_2238__delay_2237____variable_766 <= __delay_data_2238__delay_2237__delay_2236____variable_766;
      end 
      if(_mul_36_stream_oready) begin
        __delay_data_2240__delay_2239__delay_2238____variable_766 <= __delay_data_2239__delay_2238__delay_2237____variable_766;
      end 
      if(_mul_36_stream_oready) begin
        _sra_data_784 <= __muladd_data_783 >>> __delay_data_2240__delay_2239__delay_2238____variable_766;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_764 <= _cond_data_2190;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_765 <= _cond_data_1547;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_766 <= __delay_data_2874__delay_2873_plus_2241;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1525 <= _mul_36_source_start;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1526 <= _tmp_1525;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1527 <= _tmp_1526;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1528 <= _mul_36_source_start;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1529 <= _tmp_1528;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1530 <= _tmp_1529;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1531 <= _tmp_1530;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1532 <= _tmp_1531;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1533 <= _tmp_1532;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1534 <= _tmp_1533;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1535 <= _tmp_1534;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1536 <= _tmp_1535;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1537 <= _tmp_1536;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1538 <= _mul_36_source_stop;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1539 <= _tmp_1538;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1540 <= _tmp_1539;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1541 <= _tmp_1540;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1542 <= _tmp_1541;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1543 <= _tmp_1542;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1544 <= _tmp_1543;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1545 <= _tmp_1544;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1546 <= _tmp_1545;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1547 <= _tmp_1546;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1548 <= _mul_36_source_busy;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1549 <= _tmp_1548;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1550 <= _tmp_1549;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1551 <= _tmp_1550;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1552 <= _tmp_1551;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1553 <= _tmp_1552;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1554 <= _tmp_1553;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1555 <= _tmp_1554;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1556 <= _tmp_1555;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1557 <= _tmp_1556;
      end 
      if(_mul_36_stream_oready) begin
        _tmp_1558 <= _mul_36_sink_busy;
      end 
      if(!_mul_36_sink_busy && _tmp_1558) begin
        _mul_36_busy_reg <= 0;
      end 
      if(_mul_36_source_busy) begin
        _mul_36_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_36_fsm_1 = 1;
  localparam _mul_36_fsm_2 = 2;
  localparam _mul_36_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_36_fsm <= _mul_36_fsm_init;
      _mul_36_source_start <= 0;
      _mul_36_source_busy <= 0;
      _mul_36_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_36_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_36_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_36_stream_oready && _tmp_1527) begin
        _mul_36_stream_ivalid <= 1;
      end 
      if(_mul_36_stream_oready && 1'd0) begin
        _mul_36_stream_ivalid <= 0;
      end 
      case(_mul_36_fsm)
        _mul_36_fsm_init: begin
          if(_mul_36_run_flag) begin
            _mul_36_source_start <= 1;
          end 
          if(_mul_36_run_flag) begin
            _mul_36_fsm <= _mul_36_fsm_1;
          end 
        end
        _mul_36_fsm_1: begin
          if(_mul_36_source_start && _mul_36_stream_oready) begin
            _mul_36_source_start <= 0;
            _mul_36_source_busy <= 1;
          end 
          if(_mul_36_source_start && _mul_36_stream_oready) begin
            _mul_36_fsm <= _mul_36_fsm_2;
          end 
        end
        _mul_36_fsm_2: begin
          if(_mul_36_stream_oready) begin
            _mul_36_fsm <= _mul_36_fsm_3;
          end 
        end
        _mul_36_fsm_3: begin
          if(_mul_36_stream_oready && 1'd0) begin
            _mul_36_source_busy <= 0;
          end 
          if(_mul_36_stream_oready && 1'd0 && _mul_36_run_flag) begin
            _mul_36_source_start <= 1;
          end 
          if(_mul_36_stream_oready && 1'd0) begin
            _mul_36_fsm <= _mul_36_fsm_init;
          end 
          if(_mul_36_stream_oready && 1'd0 && _mul_36_run_flag) begin
            _mul_36_fsm <= _mul_36_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_37_x_source_ram_renable <= 0;
      _mul_37_x_source_fifo_deq <= 0;
      _mul_37_x_idle <= 1;
      _mul_37_y_source_ram_renable <= 0;
      _mul_37_y_source_fifo_deq <= 0;
      _mul_37_y_idle <= 1;
      _mul_37_rshift_source_ram_renable <= 0;
      _mul_37_rshift_source_fifo_deq <= 0;
      _mul_37_rshift_idle <= 1;
      _mul_37_z_sink_wenable <= 0;
      _mul_37_z_sink_fifo_enq <= 0;
      __mul_37_stream_ivalid_1 <= 0;
      __mul_37_stream_ivalid_2 <= 0;
      __mul_37_stream_ivalid_3 <= 0;
      __mul_37_stream_ivalid_4 <= 0;
      __mul_37_stream_ivalid_5 <= 0;
      __mul_37_stream_ivalid_6 <= 0;
      __mul_37_stream_ivalid_7 <= 0;
      __mul_37_stream_ivalid_8 <= 0;
      _greaterthan_data_788 <= 0;
      _minus_data_790 <= 0;
      _greatereq_data_801 <= 0;
      __delay_data_2247__variable_785 <= 0;
      __delay_data_2250__variable_786 <= 0;
      __delay_data_2253__variable_787 <= 0;
      _sll_data_792 <= 0;
      __delay_data_2244_greaterthan_788 <= 0;
      __delay_data_2245_greatereq_801 <= 0;
      __delay_data_2248__delay_2247__variable_785 <= 0;
      __delay_data_2251__delay_2250__variable_786 <= 0;
      __delay_data_2254__delay_2253__variable_787 <= 0;
      _cond_data_798 <= 0;
      __delay_data_2246__delay_2245_greatereq_801 <= 0;
      __delay_data_2249__delay_2248__delay_2247__variable_785 <= 0;
      __delay_data_2252__delay_2251__delay_2250__variable_786 <= 0;
      __delay_data_2255__delay_2254__delay_2253__variable_787 <= 0;
      __muladd_madd_odata_reg_804 <= 0;
      __delay_data_2256__delay_2255__delay_2254____variable_787 <= 0;
      __delay_data_2257__delay_2256__delay_2255____variable_787 <= 0;
      __delay_data_2258__delay_2257__delay_2256____variable_787 <= 0;
      __delay_data_2259__delay_2258__delay_2257____variable_787 <= 0;
      _sra_data_805 <= 0;
      __variable_wdata_785 <= 0;
      __variable_wdata_786 <= 0;
      __variable_wdata_787 <= 0;
      _tmp_1559 <= 0;
      _tmp_1560 <= 0;
      _tmp_1561 <= 0;
      _tmp_1562 <= 0;
      _tmp_1563 <= 0;
      _tmp_1564 <= 0;
      _tmp_1565 <= 0;
      _tmp_1566 <= 0;
      _tmp_1567 <= 0;
      _tmp_1568 <= 0;
      _tmp_1569 <= 0;
      _tmp_1570 <= 0;
      _tmp_1571 <= 0;
      _tmp_1572 <= 0;
      _tmp_1573 <= 0;
      _tmp_1574 <= 0;
      _tmp_1575 <= 0;
      _tmp_1576 <= 0;
      _tmp_1577 <= 0;
      _tmp_1578 <= 0;
      _tmp_1579 <= 0;
      _tmp_1580 <= 0;
      _tmp_1581 <= 0;
      _tmp_1582 <= 0;
      _tmp_1583 <= 0;
      _tmp_1584 <= 0;
      _tmp_1585 <= 0;
      _tmp_1586 <= 0;
      _tmp_1587 <= 0;
      _tmp_1588 <= 0;
      _tmp_1589 <= 0;
      _tmp_1590 <= 0;
      _tmp_1591 <= 0;
      _tmp_1592 <= 0;
      _mul_37_busy_reg <= 0;
    end else begin
      if(_mul_37_stream_oready) begin
        _mul_37_x_source_ram_renable <= 0;
        _mul_37_x_source_fifo_deq <= 0;
      end 
      _mul_37_x_idle <= _mul_37_x_idle;
      if(_mul_37_stream_oready) begin
        _mul_37_y_source_ram_renable <= 0;
        _mul_37_y_source_fifo_deq <= 0;
      end 
      _mul_37_y_idle <= _mul_37_y_idle;
      if(_mul_37_stream_oready) begin
        _mul_37_rshift_source_ram_renable <= 0;
        _mul_37_rshift_source_fifo_deq <= 0;
      end 
      _mul_37_rshift_idle <= _mul_37_rshift_idle;
      if(_mul_37_stream_oready) begin
        _mul_37_z_sink_wenable <= 0;
        _mul_37_z_sink_fifo_enq <= 0;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_1 <= _mul_37_stream_ivalid;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_2 <= __mul_37_stream_ivalid_1;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_3 <= __mul_37_stream_ivalid_2;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_4 <= __mul_37_stream_ivalid_3;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_5 <= __mul_37_stream_ivalid_4;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_6 <= __mul_37_stream_ivalid_5;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_7 <= __mul_37_stream_ivalid_6;
      end 
      if(_mul_37_stream_oready) begin
        __mul_37_stream_ivalid_8 <= __mul_37_stream_ivalid_7;
      end 
      if(_mul_37_stream_oready) begin
        _greaterthan_data_788 <= mul_37_rshift_data > 1'sd0;
      end 
      if(_mul_37_stream_oready) begin
        _minus_data_790 <= mul_37_rshift_data - 2'sd1;
      end 
      if(_mul_37_stream_oready) begin
        _greatereq_data_801 <= mul_37_x_data >= 1'sd0;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2247__variable_785 <= mul_37_x_data;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2250__variable_786 <= mul_37_y_data;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2253__variable_787 <= mul_37_rshift_data;
      end 
      if(_mul_37_stream_oready) begin
        _sll_data_792 <= 2'sd1 << _minus_data_790;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2244_greaterthan_788 <= _greaterthan_data_788;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2245_greatereq_801 <= _greatereq_data_801;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2248__delay_2247__variable_785 <= __delay_data_2247__variable_785;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2251__delay_2250__variable_786 <= __delay_data_2250__variable_786;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2254__delay_2253__variable_787 <= __delay_data_2253__variable_787;
      end 
      if(_mul_37_stream_oready) begin
        _cond_data_798 <= (__delay_data_2244_greaterthan_788)? _sll_data_792 : 1'sd0;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2246__delay_2245_greatereq_801 <= __delay_data_2245_greatereq_801;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2249__delay_2248__delay_2247__variable_785 <= __delay_data_2248__delay_2247__variable_785;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2252__delay_2251__delay_2250__variable_786 <= __delay_data_2251__delay_2250__variable_786;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2255__delay_2254__delay_2253__variable_787 <= __delay_data_2254__delay_2253__variable_787;
      end 
      if(_mul_37_stream_oready) begin
        __muladd_madd_odata_reg_804 <= __muladd_madd_odata_804;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2256__delay_2255__delay_2254____variable_787 <= __delay_data_2255__delay_2254__delay_2253__variable_787;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2257__delay_2256__delay_2255____variable_787 <= __delay_data_2256__delay_2255__delay_2254____variable_787;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2258__delay_2257__delay_2256____variable_787 <= __delay_data_2257__delay_2256__delay_2255____variable_787;
      end 
      if(_mul_37_stream_oready) begin
        __delay_data_2259__delay_2258__delay_2257____variable_787 <= __delay_data_2258__delay_2257__delay_2256____variable_787;
      end 
      if(_mul_37_stream_oready) begin
        _sra_data_805 <= __muladd_data_804 >>> __delay_data_2259__delay_2258__delay_2257____variable_787;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_785 <= _cond_data_2192;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_786 <= _cond_data_1549;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_787 <= __delay_data_2884__delay_2883_plus_2260;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1559 <= _mul_37_source_start;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1560 <= _tmp_1559;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1561 <= _tmp_1560;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1562 <= _mul_37_source_start;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1563 <= _tmp_1562;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1564 <= _tmp_1563;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1565 <= _tmp_1564;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1566 <= _tmp_1565;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1567 <= _tmp_1566;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1568 <= _tmp_1567;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1569 <= _tmp_1568;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1570 <= _tmp_1569;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1571 <= _tmp_1570;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1572 <= _mul_37_source_stop;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1573 <= _tmp_1572;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1574 <= _tmp_1573;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1575 <= _tmp_1574;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1576 <= _tmp_1575;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1577 <= _tmp_1576;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1578 <= _tmp_1577;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1579 <= _tmp_1578;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1580 <= _tmp_1579;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1581 <= _tmp_1580;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1582 <= _mul_37_source_busy;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1583 <= _tmp_1582;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1584 <= _tmp_1583;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1585 <= _tmp_1584;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1586 <= _tmp_1585;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1587 <= _tmp_1586;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1588 <= _tmp_1587;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1589 <= _tmp_1588;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1590 <= _tmp_1589;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1591 <= _tmp_1590;
      end 
      if(_mul_37_stream_oready) begin
        _tmp_1592 <= _mul_37_sink_busy;
      end 
      if(!_mul_37_sink_busy && _tmp_1592) begin
        _mul_37_busy_reg <= 0;
      end 
      if(_mul_37_source_busy) begin
        _mul_37_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_37_fsm_1 = 1;
  localparam _mul_37_fsm_2 = 2;
  localparam _mul_37_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_37_fsm <= _mul_37_fsm_init;
      _mul_37_source_start <= 0;
      _mul_37_source_busy <= 0;
      _mul_37_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_37_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_37_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_37_stream_oready && _tmp_1561) begin
        _mul_37_stream_ivalid <= 1;
      end 
      if(_mul_37_stream_oready && 1'd0) begin
        _mul_37_stream_ivalid <= 0;
      end 
      case(_mul_37_fsm)
        _mul_37_fsm_init: begin
          if(_mul_37_run_flag) begin
            _mul_37_source_start <= 1;
          end 
          if(_mul_37_run_flag) begin
            _mul_37_fsm <= _mul_37_fsm_1;
          end 
        end
        _mul_37_fsm_1: begin
          if(_mul_37_source_start && _mul_37_stream_oready) begin
            _mul_37_source_start <= 0;
            _mul_37_source_busy <= 1;
          end 
          if(_mul_37_source_start && _mul_37_stream_oready) begin
            _mul_37_fsm <= _mul_37_fsm_2;
          end 
        end
        _mul_37_fsm_2: begin
          if(_mul_37_stream_oready) begin
            _mul_37_fsm <= _mul_37_fsm_3;
          end 
        end
        _mul_37_fsm_3: begin
          if(_mul_37_stream_oready && 1'd0) begin
            _mul_37_source_busy <= 0;
          end 
          if(_mul_37_stream_oready && 1'd0 && _mul_37_run_flag) begin
            _mul_37_source_start <= 1;
          end 
          if(_mul_37_stream_oready && 1'd0) begin
            _mul_37_fsm <= _mul_37_fsm_init;
          end 
          if(_mul_37_stream_oready && 1'd0 && _mul_37_run_flag) begin
            _mul_37_fsm <= _mul_37_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_38_x_source_ram_renable <= 0;
      _mul_38_x_source_fifo_deq <= 0;
      _mul_38_x_idle <= 1;
      _mul_38_y_source_ram_renable <= 0;
      _mul_38_y_source_fifo_deq <= 0;
      _mul_38_y_idle <= 1;
      _mul_38_rshift_source_ram_renable <= 0;
      _mul_38_rshift_source_fifo_deq <= 0;
      _mul_38_rshift_idle <= 1;
      _mul_38_z_sink_wenable <= 0;
      _mul_38_z_sink_fifo_enq <= 0;
      __mul_38_stream_ivalid_1 <= 0;
      __mul_38_stream_ivalid_2 <= 0;
      __mul_38_stream_ivalid_3 <= 0;
      __mul_38_stream_ivalid_4 <= 0;
      __mul_38_stream_ivalid_5 <= 0;
      __mul_38_stream_ivalid_6 <= 0;
      __mul_38_stream_ivalid_7 <= 0;
      __mul_38_stream_ivalid_8 <= 0;
      _greaterthan_data_809 <= 0;
      _minus_data_811 <= 0;
      _greatereq_data_822 <= 0;
      __delay_data_2266__variable_806 <= 0;
      __delay_data_2269__variable_807 <= 0;
      __delay_data_2272__variable_808 <= 0;
      _sll_data_813 <= 0;
      __delay_data_2263_greaterthan_809 <= 0;
      __delay_data_2264_greatereq_822 <= 0;
      __delay_data_2267__delay_2266__variable_806 <= 0;
      __delay_data_2270__delay_2269__variable_807 <= 0;
      __delay_data_2273__delay_2272__variable_808 <= 0;
      _cond_data_819 <= 0;
      __delay_data_2265__delay_2264_greatereq_822 <= 0;
      __delay_data_2268__delay_2267__delay_2266__variable_806 <= 0;
      __delay_data_2271__delay_2270__delay_2269__variable_807 <= 0;
      __delay_data_2274__delay_2273__delay_2272__variable_808 <= 0;
      __muladd_madd_odata_reg_825 <= 0;
      __delay_data_2275__delay_2274__delay_2273____variable_808 <= 0;
      __delay_data_2276__delay_2275__delay_2274____variable_808 <= 0;
      __delay_data_2277__delay_2276__delay_2275____variable_808 <= 0;
      __delay_data_2278__delay_2277__delay_2276____variable_808 <= 0;
      _sra_data_826 <= 0;
      __variable_wdata_806 <= 0;
      __variable_wdata_807 <= 0;
      __variable_wdata_808 <= 0;
      _tmp_1593 <= 0;
      _tmp_1594 <= 0;
      _tmp_1595 <= 0;
      _tmp_1596 <= 0;
      _tmp_1597 <= 0;
      _tmp_1598 <= 0;
      _tmp_1599 <= 0;
      _tmp_1600 <= 0;
      _tmp_1601 <= 0;
      _tmp_1602 <= 0;
      _tmp_1603 <= 0;
      _tmp_1604 <= 0;
      _tmp_1605 <= 0;
      _tmp_1606 <= 0;
      _tmp_1607 <= 0;
      _tmp_1608 <= 0;
      _tmp_1609 <= 0;
      _tmp_1610 <= 0;
      _tmp_1611 <= 0;
      _tmp_1612 <= 0;
      _tmp_1613 <= 0;
      _tmp_1614 <= 0;
      _tmp_1615 <= 0;
      _tmp_1616 <= 0;
      _tmp_1617 <= 0;
      _tmp_1618 <= 0;
      _tmp_1619 <= 0;
      _tmp_1620 <= 0;
      _tmp_1621 <= 0;
      _tmp_1622 <= 0;
      _tmp_1623 <= 0;
      _tmp_1624 <= 0;
      _tmp_1625 <= 0;
      _tmp_1626 <= 0;
      _mul_38_busy_reg <= 0;
    end else begin
      if(_mul_38_stream_oready) begin
        _mul_38_x_source_ram_renable <= 0;
        _mul_38_x_source_fifo_deq <= 0;
      end 
      _mul_38_x_idle <= _mul_38_x_idle;
      if(_mul_38_stream_oready) begin
        _mul_38_y_source_ram_renable <= 0;
        _mul_38_y_source_fifo_deq <= 0;
      end 
      _mul_38_y_idle <= _mul_38_y_idle;
      if(_mul_38_stream_oready) begin
        _mul_38_rshift_source_ram_renable <= 0;
        _mul_38_rshift_source_fifo_deq <= 0;
      end 
      _mul_38_rshift_idle <= _mul_38_rshift_idle;
      if(_mul_38_stream_oready) begin
        _mul_38_z_sink_wenable <= 0;
        _mul_38_z_sink_fifo_enq <= 0;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_1 <= _mul_38_stream_ivalid;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_2 <= __mul_38_stream_ivalid_1;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_3 <= __mul_38_stream_ivalid_2;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_4 <= __mul_38_stream_ivalid_3;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_5 <= __mul_38_stream_ivalid_4;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_6 <= __mul_38_stream_ivalid_5;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_7 <= __mul_38_stream_ivalid_6;
      end 
      if(_mul_38_stream_oready) begin
        __mul_38_stream_ivalid_8 <= __mul_38_stream_ivalid_7;
      end 
      if(_mul_38_stream_oready) begin
        _greaterthan_data_809 <= mul_38_rshift_data > 1'sd0;
      end 
      if(_mul_38_stream_oready) begin
        _minus_data_811 <= mul_38_rshift_data - 2'sd1;
      end 
      if(_mul_38_stream_oready) begin
        _greatereq_data_822 <= mul_38_x_data >= 1'sd0;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2266__variable_806 <= mul_38_x_data;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2269__variable_807 <= mul_38_y_data;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2272__variable_808 <= mul_38_rshift_data;
      end 
      if(_mul_38_stream_oready) begin
        _sll_data_813 <= 2'sd1 << _minus_data_811;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2263_greaterthan_809 <= _greaterthan_data_809;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2264_greatereq_822 <= _greatereq_data_822;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2267__delay_2266__variable_806 <= __delay_data_2266__variable_806;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2270__delay_2269__variable_807 <= __delay_data_2269__variable_807;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2273__delay_2272__variable_808 <= __delay_data_2272__variable_808;
      end 
      if(_mul_38_stream_oready) begin
        _cond_data_819 <= (__delay_data_2263_greaterthan_809)? _sll_data_813 : 1'sd0;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2265__delay_2264_greatereq_822 <= __delay_data_2264_greatereq_822;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2268__delay_2267__delay_2266__variable_806 <= __delay_data_2267__delay_2266__variable_806;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2271__delay_2270__delay_2269__variable_807 <= __delay_data_2270__delay_2269__variable_807;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2274__delay_2273__delay_2272__variable_808 <= __delay_data_2273__delay_2272__variable_808;
      end 
      if(_mul_38_stream_oready) begin
        __muladd_madd_odata_reg_825 <= __muladd_madd_odata_825;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2275__delay_2274__delay_2273____variable_808 <= __delay_data_2274__delay_2273__delay_2272__variable_808;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2276__delay_2275__delay_2274____variable_808 <= __delay_data_2275__delay_2274__delay_2273____variable_808;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2277__delay_2276__delay_2275____variable_808 <= __delay_data_2276__delay_2275__delay_2274____variable_808;
      end 
      if(_mul_38_stream_oready) begin
        __delay_data_2278__delay_2277__delay_2276____variable_808 <= __delay_data_2277__delay_2276__delay_2275____variable_808;
      end 
      if(_mul_38_stream_oready) begin
        _sra_data_826 <= __muladd_data_825 >>> __delay_data_2278__delay_2277__delay_2276____variable_808;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_806 <= _cond_data_2194;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_807 <= _cond_data_1551;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_808 <= __delay_data_2894__delay_2893_plus_2279;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1593 <= _mul_38_source_start;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1594 <= _tmp_1593;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1595 <= _tmp_1594;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1596 <= _mul_38_source_start;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1597 <= _tmp_1596;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1598 <= _tmp_1597;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1599 <= _tmp_1598;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1600 <= _tmp_1599;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1601 <= _tmp_1600;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1602 <= _tmp_1601;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1603 <= _tmp_1602;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1604 <= _tmp_1603;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1605 <= _tmp_1604;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1606 <= _mul_38_source_stop;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1607 <= _tmp_1606;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1608 <= _tmp_1607;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1609 <= _tmp_1608;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1610 <= _tmp_1609;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1611 <= _tmp_1610;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1612 <= _tmp_1611;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1613 <= _tmp_1612;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1614 <= _tmp_1613;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1615 <= _tmp_1614;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1616 <= _mul_38_source_busy;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1617 <= _tmp_1616;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1618 <= _tmp_1617;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1619 <= _tmp_1618;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1620 <= _tmp_1619;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1621 <= _tmp_1620;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1622 <= _tmp_1621;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1623 <= _tmp_1622;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1624 <= _tmp_1623;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1625 <= _tmp_1624;
      end 
      if(_mul_38_stream_oready) begin
        _tmp_1626 <= _mul_38_sink_busy;
      end 
      if(!_mul_38_sink_busy && _tmp_1626) begin
        _mul_38_busy_reg <= 0;
      end 
      if(_mul_38_source_busy) begin
        _mul_38_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_38_fsm_1 = 1;
  localparam _mul_38_fsm_2 = 2;
  localparam _mul_38_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_38_fsm <= _mul_38_fsm_init;
      _mul_38_source_start <= 0;
      _mul_38_source_busy <= 0;
      _mul_38_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_38_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_38_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_38_stream_oready && _tmp_1595) begin
        _mul_38_stream_ivalid <= 1;
      end 
      if(_mul_38_stream_oready && 1'd0) begin
        _mul_38_stream_ivalid <= 0;
      end 
      case(_mul_38_fsm)
        _mul_38_fsm_init: begin
          if(_mul_38_run_flag) begin
            _mul_38_source_start <= 1;
          end 
          if(_mul_38_run_flag) begin
            _mul_38_fsm <= _mul_38_fsm_1;
          end 
        end
        _mul_38_fsm_1: begin
          if(_mul_38_source_start && _mul_38_stream_oready) begin
            _mul_38_source_start <= 0;
            _mul_38_source_busy <= 1;
          end 
          if(_mul_38_source_start && _mul_38_stream_oready) begin
            _mul_38_fsm <= _mul_38_fsm_2;
          end 
        end
        _mul_38_fsm_2: begin
          if(_mul_38_stream_oready) begin
            _mul_38_fsm <= _mul_38_fsm_3;
          end 
        end
        _mul_38_fsm_3: begin
          if(_mul_38_stream_oready && 1'd0) begin
            _mul_38_source_busy <= 0;
          end 
          if(_mul_38_stream_oready && 1'd0 && _mul_38_run_flag) begin
            _mul_38_source_start <= 1;
          end 
          if(_mul_38_stream_oready && 1'd0) begin
            _mul_38_fsm <= _mul_38_fsm_init;
          end 
          if(_mul_38_stream_oready && 1'd0 && _mul_38_run_flag) begin
            _mul_38_fsm <= _mul_38_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_39_x_source_ram_renable <= 0;
      _mul_39_x_source_fifo_deq <= 0;
      _mul_39_x_idle <= 1;
      _mul_39_y_source_ram_renable <= 0;
      _mul_39_y_source_fifo_deq <= 0;
      _mul_39_y_idle <= 1;
      _mul_39_rshift_source_ram_renable <= 0;
      _mul_39_rshift_source_fifo_deq <= 0;
      _mul_39_rshift_idle <= 1;
      _mul_39_z_sink_wenable <= 0;
      _mul_39_z_sink_fifo_enq <= 0;
      __mul_39_stream_ivalid_1 <= 0;
      __mul_39_stream_ivalid_2 <= 0;
      __mul_39_stream_ivalid_3 <= 0;
      __mul_39_stream_ivalid_4 <= 0;
      __mul_39_stream_ivalid_5 <= 0;
      __mul_39_stream_ivalid_6 <= 0;
      __mul_39_stream_ivalid_7 <= 0;
      __mul_39_stream_ivalid_8 <= 0;
      _greaterthan_data_830 <= 0;
      _minus_data_832 <= 0;
      _greatereq_data_843 <= 0;
      __delay_data_2285__variable_827 <= 0;
      __delay_data_2288__variable_828 <= 0;
      __delay_data_2291__variable_829 <= 0;
      _sll_data_834 <= 0;
      __delay_data_2282_greaterthan_830 <= 0;
      __delay_data_2283_greatereq_843 <= 0;
      __delay_data_2286__delay_2285__variable_827 <= 0;
      __delay_data_2289__delay_2288__variable_828 <= 0;
      __delay_data_2292__delay_2291__variable_829 <= 0;
      _cond_data_840 <= 0;
      __delay_data_2284__delay_2283_greatereq_843 <= 0;
      __delay_data_2287__delay_2286__delay_2285__variable_827 <= 0;
      __delay_data_2290__delay_2289__delay_2288__variable_828 <= 0;
      __delay_data_2293__delay_2292__delay_2291__variable_829 <= 0;
      __muladd_madd_odata_reg_846 <= 0;
      __delay_data_2294__delay_2293__delay_2292____variable_829 <= 0;
      __delay_data_2295__delay_2294__delay_2293____variable_829 <= 0;
      __delay_data_2296__delay_2295__delay_2294____variable_829 <= 0;
      __delay_data_2297__delay_2296__delay_2295____variable_829 <= 0;
      _sra_data_847 <= 0;
      __variable_wdata_827 <= 0;
      __variable_wdata_828 <= 0;
      __variable_wdata_829 <= 0;
      _tmp_1627 <= 0;
      _tmp_1628 <= 0;
      _tmp_1629 <= 0;
      _tmp_1630 <= 0;
      _tmp_1631 <= 0;
      _tmp_1632 <= 0;
      _tmp_1633 <= 0;
      _tmp_1634 <= 0;
      _tmp_1635 <= 0;
      _tmp_1636 <= 0;
      _tmp_1637 <= 0;
      _tmp_1638 <= 0;
      _tmp_1639 <= 0;
      _tmp_1640 <= 0;
      _tmp_1641 <= 0;
      _tmp_1642 <= 0;
      _tmp_1643 <= 0;
      _tmp_1644 <= 0;
      _tmp_1645 <= 0;
      _tmp_1646 <= 0;
      _tmp_1647 <= 0;
      _tmp_1648 <= 0;
      _tmp_1649 <= 0;
      _tmp_1650 <= 0;
      _tmp_1651 <= 0;
      _tmp_1652 <= 0;
      _tmp_1653 <= 0;
      _tmp_1654 <= 0;
      _tmp_1655 <= 0;
      _tmp_1656 <= 0;
      _tmp_1657 <= 0;
      _tmp_1658 <= 0;
      _tmp_1659 <= 0;
      _tmp_1660 <= 0;
      _mul_39_busy_reg <= 0;
    end else begin
      if(_mul_39_stream_oready) begin
        _mul_39_x_source_ram_renable <= 0;
        _mul_39_x_source_fifo_deq <= 0;
      end 
      _mul_39_x_idle <= _mul_39_x_idle;
      if(_mul_39_stream_oready) begin
        _mul_39_y_source_ram_renable <= 0;
        _mul_39_y_source_fifo_deq <= 0;
      end 
      _mul_39_y_idle <= _mul_39_y_idle;
      if(_mul_39_stream_oready) begin
        _mul_39_rshift_source_ram_renable <= 0;
        _mul_39_rshift_source_fifo_deq <= 0;
      end 
      _mul_39_rshift_idle <= _mul_39_rshift_idle;
      if(_mul_39_stream_oready) begin
        _mul_39_z_sink_wenable <= 0;
        _mul_39_z_sink_fifo_enq <= 0;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_1 <= _mul_39_stream_ivalid;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_2 <= __mul_39_stream_ivalid_1;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_3 <= __mul_39_stream_ivalid_2;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_4 <= __mul_39_stream_ivalid_3;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_5 <= __mul_39_stream_ivalid_4;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_6 <= __mul_39_stream_ivalid_5;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_7 <= __mul_39_stream_ivalid_6;
      end 
      if(_mul_39_stream_oready) begin
        __mul_39_stream_ivalid_8 <= __mul_39_stream_ivalid_7;
      end 
      if(_mul_39_stream_oready) begin
        _greaterthan_data_830 <= mul_39_rshift_data > 1'sd0;
      end 
      if(_mul_39_stream_oready) begin
        _minus_data_832 <= mul_39_rshift_data - 2'sd1;
      end 
      if(_mul_39_stream_oready) begin
        _greatereq_data_843 <= mul_39_x_data >= 1'sd0;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2285__variable_827 <= mul_39_x_data;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2288__variable_828 <= mul_39_y_data;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2291__variable_829 <= mul_39_rshift_data;
      end 
      if(_mul_39_stream_oready) begin
        _sll_data_834 <= 2'sd1 << _minus_data_832;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2282_greaterthan_830 <= _greaterthan_data_830;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2283_greatereq_843 <= _greatereq_data_843;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2286__delay_2285__variable_827 <= __delay_data_2285__variable_827;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2289__delay_2288__variable_828 <= __delay_data_2288__variable_828;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2292__delay_2291__variable_829 <= __delay_data_2291__variable_829;
      end 
      if(_mul_39_stream_oready) begin
        _cond_data_840 <= (__delay_data_2282_greaterthan_830)? _sll_data_834 : 1'sd0;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2284__delay_2283_greatereq_843 <= __delay_data_2283_greatereq_843;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2287__delay_2286__delay_2285__variable_827 <= __delay_data_2286__delay_2285__variable_827;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2290__delay_2289__delay_2288__variable_828 <= __delay_data_2289__delay_2288__variable_828;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2293__delay_2292__delay_2291__variable_829 <= __delay_data_2292__delay_2291__variable_829;
      end 
      if(_mul_39_stream_oready) begin
        __muladd_madd_odata_reg_846 <= __muladd_madd_odata_846;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2294__delay_2293__delay_2292____variable_829 <= __delay_data_2293__delay_2292__delay_2291__variable_829;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2295__delay_2294__delay_2293____variable_829 <= __delay_data_2294__delay_2293__delay_2292____variable_829;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2296__delay_2295__delay_2294____variable_829 <= __delay_data_2295__delay_2294__delay_2293____variable_829;
      end 
      if(_mul_39_stream_oready) begin
        __delay_data_2297__delay_2296__delay_2295____variable_829 <= __delay_data_2296__delay_2295__delay_2294____variable_829;
      end 
      if(_mul_39_stream_oready) begin
        _sra_data_847 <= __muladd_data_846 >>> __delay_data_2297__delay_2296__delay_2295____variable_829;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_827 <= _cond_data_2196;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_828 <= _cond_data_1553;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_829 <= __delay_data_2904__delay_2903_plus_2298;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1627 <= _mul_39_source_start;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1628 <= _tmp_1627;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1629 <= _tmp_1628;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1630 <= _mul_39_source_start;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1631 <= _tmp_1630;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1632 <= _tmp_1631;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1633 <= _tmp_1632;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1634 <= _tmp_1633;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1635 <= _tmp_1634;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1636 <= _tmp_1635;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1637 <= _tmp_1636;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1638 <= _tmp_1637;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1639 <= _tmp_1638;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1640 <= _mul_39_source_stop;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1641 <= _tmp_1640;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1642 <= _tmp_1641;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1643 <= _tmp_1642;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1644 <= _tmp_1643;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1645 <= _tmp_1644;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1646 <= _tmp_1645;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1647 <= _tmp_1646;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1648 <= _tmp_1647;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1649 <= _tmp_1648;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1650 <= _mul_39_source_busy;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1651 <= _tmp_1650;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1652 <= _tmp_1651;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1653 <= _tmp_1652;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1654 <= _tmp_1653;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1655 <= _tmp_1654;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1656 <= _tmp_1655;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1657 <= _tmp_1656;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1658 <= _tmp_1657;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1659 <= _tmp_1658;
      end 
      if(_mul_39_stream_oready) begin
        _tmp_1660 <= _mul_39_sink_busy;
      end 
      if(!_mul_39_sink_busy && _tmp_1660) begin
        _mul_39_busy_reg <= 0;
      end 
      if(_mul_39_source_busy) begin
        _mul_39_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_39_fsm_1 = 1;
  localparam _mul_39_fsm_2 = 2;
  localparam _mul_39_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_39_fsm <= _mul_39_fsm_init;
      _mul_39_source_start <= 0;
      _mul_39_source_busy <= 0;
      _mul_39_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_39_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_39_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_39_stream_oready && _tmp_1629) begin
        _mul_39_stream_ivalid <= 1;
      end 
      if(_mul_39_stream_oready && 1'd0) begin
        _mul_39_stream_ivalid <= 0;
      end 
      case(_mul_39_fsm)
        _mul_39_fsm_init: begin
          if(_mul_39_run_flag) begin
            _mul_39_source_start <= 1;
          end 
          if(_mul_39_run_flag) begin
            _mul_39_fsm <= _mul_39_fsm_1;
          end 
        end
        _mul_39_fsm_1: begin
          if(_mul_39_source_start && _mul_39_stream_oready) begin
            _mul_39_source_start <= 0;
            _mul_39_source_busy <= 1;
          end 
          if(_mul_39_source_start && _mul_39_stream_oready) begin
            _mul_39_fsm <= _mul_39_fsm_2;
          end 
        end
        _mul_39_fsm_2: begin
          if(_mul_39_stream_oready) begin
            _mul_39_fsm <= _mul_39_fsm_3;
          end 
        end
        _mul_39_fsm_3: begin
          if(_mul_39_stream_oready && 1'd0) begin
            _mul_39_source_busy <= 0;
          end 
          if(_mul_39_stream_oready && 1'd0 && _mul_39_run_flag) begin
            _mul_39_source_start <= 1;
          end 
          if(_mul_39_stream_oready && 1'd0) begin
            _mul_39_fsm <= _mul_39_fsm_init;
          end 
          if(_mul_39_stream_oready && 1'd0 && _mul_39_run_flag) begin
            _mul_39_fsm <= _mul_39_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_40_x_source_ram_renable <= 0;
      _mul_40_x_source_fifo_deq <= 0;
      _mul_40_x_idle <= 1;
      _mul_40_y_source_ram_renable <= 0;
      _mul_40_y_source_fifo_deq <= 0;
      _mul_40_y_idle <= 1;
      _mul_40_rshift_source_ram_renable <= 0;
      _mul_40_rshift_source_fifo_deq <= 0;
      _mul_40_rshift_idle <= 1;
      _mul_40_z_sink_wenable <= 0;
      _mul_40_z_sink_fifo_enq <= 0;
      __mul_40_stream_ivalid_1 <= 0;
      __mul_40_stream_ivalid_2 <= 0;
      __mul_40_stream_ivalid_3 <= 0;
      __mul_40_stream_ivalid_4 <= 0;
      __mul_40_stream_ivalid_5 <= 0;
      __mul_40_stream_ivalid_6 <= 0;
      __mul_40_stream_ivalid_7 <= 0;
      __mul_40_stream_ivalid_8 <= 0;
      _greaterthan_data_851 <= 0;
      _minus_data_853 <= 0;
      _greatereq_data_864 <= 0;
      __delay_data_2304__variable_848 <= 0;
      __delay_data_2307__variable_849 <= 0;
      __delay_data_2310__variable_850 <= 0;
      _sll_data_855 <= 0;
      __delay_data_2301_greaterthan_851 <= 0;
      __delay_data_2302_greatereq_864 <= 0;
      __delay_data_2305__delay_2304__variable_848 <= 0;
      __delay_data_2308__delay_2307__variable_849 <= 0;
      __delay_data_2311__delay_2310__variable_850 <= 0;
      _cond_data_861 <= 0;
      __delay_data_2303__delay_2302_greatereq_864 <= 0;
      __delay_data_2306__delay_2305__delay_2304__variable_848 <= 0;
      __delay_data_2309__delay_2308__delay_2307__variable_849 <= 0;
      __delay_data_2312__delay_2311__delay_2310__variable_850 <= 0;
      __muladd_madd_odata_reg_867 <= 0;
      __delay_data_2313__delay_2312__delay_2311____variable_850 <= 0;
      __delay_data_2314__delay_2313__delay_2312____variable_850 <= 0;
      __delay_data_2315__delay_2314__delay_2313____variable_850 <= 0;
      __delay_data_2316__delay_2315__delay_2314____variable_850 <= 0;
      _sra_data_868 <= 0;
      __variable_wdata_848 <= 0;
      __variable_wdata_849 <= 0;
      __variable_wdata_850 <= 0;
      _tmp_1661 <= 0;
      _tmp_1662 <= 0;
      _tmp_1663 <= 0;
      _tmp_1664 <= 0;
      _tmp_1665 <= 0;
      _tmp_1666 <= 0;
      _tmp_1667 <= 0;
      _tmp_1668 <= 0;
      _tmp_1669 <= 0;
      _tmp_1670 <= 0;
      _tmp_1671 <= 0;
      _tmp_1672 <= 0;
      _tmp_1673 <= 0;
      _tmp_1674 <= 0;
      _tmp_1675 <= 0;
      _tmp_1676 <= 0;
      _tmp_1677 <= 0;
      _tmp_1678 <= 0;
      _tmp_1679 <= 0;
      _tmp_1680 <= 0;
      _tmp_1681 <= 0;
      _tmp_1682 <= 0;
      _tmp_1683 <= 0;
      _tmp_1684 <= 0;
      _tmp_1685 <= 0;
      _tmp_1686 <= 0;
      _tmp_1687 <= 0;
      _tmp_1688 <= 0;
      _tmp_1689 <= 0;
      _tmp_1690 <= 0;
      _tmp_1691 <= 0;
      _tmp_1692 <= 0;
      _tmp_1693 <= 0;
      _tmp_1694 <= 0;
      _mul_40_busy_reg <= 0;
    end else begin
      if(_mul_40_stream_oready) begin
        _mul_40_x_source_ram_renable <= 0;
        _mul_40_x_source_fifo_deq <= 0;
      end 
      _mul_40_x_idle <= _mul_40_x_idle;
      if(_mul_40_stream_oready) begin
        _mul_40_y_source_ram_renable <= 0;
        _mul_40_y_source_fifo_deq <= 0;
      end 
      _mul_40_y_idle <= _mul_40_y_idle;
      if(_mul_40_stream_oready) begin
        _mul_40_rshift_source_ram_renable <= 0;
        _mul_40_rshift_source_fifo_deq <= 0;
      end 
      _mul_40_rshift_idle <= _mul_40_rshift_idle;
      if(_mul_40_stream_oready) begin
        _mul_40_z_sink_wenable <= 0;
        _mul_40_z_sink_fifo_enq <= 0;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_1 <= _mul_40_stream_ivalid;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_2 <= __mul_40_stream_ivalid_1;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_3 <= __mul_40_stream_ivalid_2;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_4 <= __mul_40_stream_ivalid_3;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_5 <= __mul_40_stream_ivalid_4;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_6 <= __mul_40_stream_ivalid_5;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_7 <= __mul_40_stream_ivalid_6;
      end 
      if(_mul_40_stream_oready) begin
        __mul_40_stream_ivalid_8 <= __mul_40_stream_ivalid_7;
      end 
      if(_mul_40_stream_oready) begin
        _greaterthan_data_851 <= mul_40_rshift_data > 1'sd0;
      end 
      if(_mul_40_stream_oready) begin
        _minus_data_853 <= mul_40_rshift_data - 2'sd1;
      end 
      if(_mul_40_stream_oready) begin
        _greatereq_data_864 <= mul_40_x_data >= 1'sd0;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2304__variable_848 <= mul_40_x_data;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2307__variable_849 <= mul_40_y_data;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2310__variable_850 <= mul_40_rshift_data;
      end 
      if(_mul_40_stream_oready) begin
        _sll_data_855 <= 2'sd1 << _minus_data_853;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2301_greaterthan_851 <= _greaterthan_data_851;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2302_greatereq_864 <= _greatereq_data_864;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2305__delay_2304__variable_848 <= __delay_data_2304__variable_848;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2308__delay_2307__variable_849 <= __delay_data_2307__variable_849;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2311__delay_2310__variable_850 <= __delay_data_2310__variable_850;
      end 
      if(_mul_40_stream_oready) begin
        _cond_data_861 <= (__delay_data_2301_greaterthan_851)? _sll_data_855 : 1'sd0;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2303__delay_2302_greatereq_864 <= __delay_data_2302_greatereq_864;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2306__delay_2305__delay_2304__variable_848 <= __delay_data_2305__delay_2304__variable_848;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2309__delay_2308__delay_2307__variable_849 <= __delay_data_2308__delay_2307__variable_849;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2312__delay_2311__delay_2310__variable_850 <= __delay_data_2311__delay_2310__variable_850;
      end 
      if(_mul_40_stream_oready) begin
        __muladd_madd_odata_reg_867 <= __muladd_madd_odata_867;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2313__delay_2312__delay_2311____variable_850 <= __delay_data_2312__delay_2311__delay_2310__variable_850;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2314__delay_2313__delay_2312____variable_850 <= __delay_data_2313__delay_2312__delay_2311____variable_850;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2315__delay_2314__delay_2313____variable_850 <= __delay_data_2314__delay_2313__delay_2312____variable_850;
      end 
      if(_mul_40_stream_oready) begin
        __delay_data_2316__delay_2315__delay_2314____variable_850 <= __delay_data_2315__delay_2314__delay_2313____variable_850;
      end 
      if(_mul_40_stream_oready) begin
        _sra_data_868 <= __muladd_data_867 >>> __delay_data_2316__delay_2315__delay_2314____variable_850;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_848 <= _cond_data_2198;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_849 <= _cond_data_1555;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_850 <= __delay_data_2914__delay_2913_plus_2317;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1661 <= _mul_40_source_start;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1662 <= _tmp_1661;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1663 <= _tmp_1662;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1664 <= _mul_40_source_start;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1665 <= _tmp_1664;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1666 <= _tmp_1665;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1667 <= _tmp_1666;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1668 <= _tmp_1667;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1669 <= _tmp_1668;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1670 <= _tmp_1669;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1671 <= _tmp_1670;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1672 <= _tmp_1671;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1673 <= _tmp_1672;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1674 <= _mul_40_source_stop;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1675 <= _tmp_1674;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1676 <= _tmp_1675;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1677 <= _tmp_1676;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1678 <= _tmp_1677;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1679 <= _tmp_1678;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1680 <= _tmp_1679;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1681 <= _tmp_1680;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1682 <= _tmp_1681;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1683 <= _tmp_1682;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1684 <= _mul_40_source_busy;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1685 <= _tmp_1684;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1686 <= _tmp_1685;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1687 <= _tmp_1686;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1688 <= _tmp_1687;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1689 <= _tmp_1688;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1690 <= _tmp_1689;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1691 <= _tmp_1690;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1692 <= _tmp_1691;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1693 <= _tmp_1692;
      end 
      if(_mul_40_stream_oready) begin
        _tmp_1694 <= _mul_40_sink_busy;
      end 
      if(!_mul_40_sink_busy && _tmp_1694) begin
        _mul_40_busy_reg <= 0;
      end 
      if(_mul_40_source_busy) begin
        _mul_40_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_40_fsm_1 = 1;
  localparam _mul_40_fsm_2 = 2;
  localparam _mul_40_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_40_fsm <= _mul_40_fsm_init;
      _mul_40_source_start <= 0;
      _mul_40_source_busy <= 0;
      _mul_40_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_40_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_40_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_40_stream_oready && _tmp_1663) begin
        _mul_40_stream_ivalid <= 1;
      end 
      if(_mul_40_stream_oready && 1'd0) begin
        _mul_40_stream_ivalid <= 0;
      end 
      case(_mul_40_fsm)
        _mul_40_fsm_init: begin
          if(_mul_40_run_flag) begin
            _mul_40_source_start <= 1;
          end 
          if(_mul_40_run_flag) begin
            _mul_40_fsm <= _mul_40_fsm_1;
          end 
        end
        _mul_40_fsm_1: begin
          if(_mul_40_source_start && _mul_40_stream_oready) begin
            _mul_40_source_start <= 0;
            _mul_40_source_busy <= 1;
          end 
          if(_mul_40_source_start && _mul_40_stream_oready) begin
            _mul_40_fsm <= _mul_40_fsm_2;
          end 
        end
        _mul_40_fsm_2: begin
          if(_mul_40_stream_oready) begin
            _mul_40_fsm <= _mul_40_fsm_3;
          end 
        end
        _mul_40_fsm_3: begin
          if(_mul_40_stream_oready && 1'd0) begin
            _mul_40_source_busy <= 0;
          end 
          if(_mul_40_stream_oready && 1'd0 && _mul_40_run_flag) begin
            _mul_40_source_start <= 1;
          end 
          if(_mul_40_stream_oready && 1'd0) begin
            _mul_40_fsm <= _mul_40_fsm_init;
          end 
          if(_mul_40_stream_oready && 1'd0 && _mul_40_run_flag) begin
            _mul_40_fsm <= _mul_40_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_41_x_source_ram_renable <= 0;
      _mul_41_x_source_fifo_deq <= 0;
      _mul_41_x_idle <= 1;
      _mul_41_y_source_ram_renable <= 0;
      _mul_41_y_source_fifo_deq <= 0;
      _mul_41_y_idle <= 1;
      _mul_41_rshift_source_ram_renable <= 0;
      _mul_41_rshift_source_fifo_deq <= 0;
      _mul_41_rshift_idle <= 1;
      _mul_41_z_sink_wenable <= 0;
      _mul_41_z_sink_fifo_enq <= 0;
      __mul_41_stream_ivalid_1 <= 0;
      __mul_41_stream_ivalid_2 <= 0;
      __mul_41_stream_ivalid_3 <= 0;
      __mul_41_stream_ivalid_4 <= 0;
      __mul_41_stream_ivalid_5 <= 0;
      __mul_41_stream_ivalid_6 <= 0;
      __mul_41_stream_ivalid_7 <= 0;
      __mul_41_stream_ivalid_8 <= 0;
      _greaterthan_data_872 <= 0;
      _minus_data_874 <= 0;
      _greatereq_data_885 <= 0;
      __delay_data_2323__variable_869 <= 0;
      __delay_data_2326__variable_870 <= 0;
      __delay_data_2329__variable_871 <= 0;
      _sll_data_876 <= 0;
      __delay_data_2320_greaterthan_872 <= 0;
      __delay_data_2321_greatereq_885 <= 0;
      __delay_data_2324__delay_2323__variable_869 <= 0;
      __delay_data_2327__delay_2326__variable_870 <= 0;
      __delay_data_2330__delay_2329__variable_871 <= 0;
      _cond_data_882 <= 0;
      __delay_data_2322__delay_2321_greatereq_885 <= 0;
      __delay_data_2325__delay_2324__delay_2323__variable_869 <= 0;
      __delay_data_2328__delay_2327__delay_2326__variable_870 <= 0;
      __delay_data_2331__delay_2330__delay_2329__variable_871 <= 0;
      __muladd_madd_odata_reg_888 <= 0;
      __delay_data_2332__delay_2331__delay_2330____variable_871 <= 0;
      __delay_data_2333__delay_2332__delay_2331____variable_871 <= 0;
      __delay_data_2334__delay_2333__delay_2332____variable_871 <= 0;
      __delay_data_2335__delay_2334__delay_2333____variable_871 <= 0;
      _sra_data_889 <= 0;
      __variable_wdata_869 <= 0;
      __variable_wdata_870 <= 0;
      __variable_wdata_871 <= 0;
      _tmp_1695 <= 0;
      _tmp_1696 <= 0;
      _tmp_1697 <= 0;
      _tmp_1698 <= 0;
      _tmp_1699 <= 0;
      _tmp_1700 <= 0;
      _tmp_1701 <= 0;
      _tmp_1702 <= 0;
      _tmp_1703 <= 0;
      _tmp_1704 <= 0;
      _tmp_1705 <= 0;
      _tmp_1706 <= 0;
      _tmp_1707 <= 0;
      _tmp_1708 <= 0;
      _tmp_1709 <= 0;
      _tmp_1710 <= 0;
      _tmp_1711 <= 0;
      _tmp_1712 <= 0;
      _tmp_1713 <= 0;
      _tmp_1714 <= 0;
      _tmp_1715 <= 0;
      _tmp_1716 <= 0;
      _tmp_1717 <= 0;
      _tmp_1718 <= 0;
      _tmp_1719 <= 0;
      _tmp_1720 <= 0;
      _tmp_1721 <= 0;
      _tmp_1722 <= 0;
      _tmp_1723 <= 0;
      _tmp_1724 <= 0;
      _tmp_1725 <= 0;
      _tmp_1726 <= 0;
      _tmp_1727 <= 0;
      _tmp_1728 <= 0;
      _mul_41_busy_reg <= 0;
    end else begin
      if(_mul_41_stream_oready) begin
        _mul_41_x_source_ram_renable <= 0;
        _mul_41_x_source_fifo_deq <= 0;
      end 
      _mul_41_x_idle <= _mul_41_x_idle;
      if(_mul_41_stream_oready) begin
        _mul_41_y_source_ram_renable <= 0;
        _mul_41_y_source_fifo_deq <= 0;
      end 
      _mul_41_y_idle <= _mul_41_y_idle;
      if(_mul_41_stream_oready) begin
        _mul_41_rshift_source_ram_renable <= 0;
        _mul_41_rshift_source_fifo_deq <= 0;
      end 
      _mul_41_rshift_idle <= _mul_41_rshift_idle;
      if(_mul_41_stream_oready) begin
        _mul_41_z_sink_wenable <= 0;
        _mul_41_z_sink_fifo_enq <= 0;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_1 <= _mul_41_stream_ivalid;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_2 <= __mul_41_stream_ivalid_1;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_3 <= __mul_41_stream_ivalid_2;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_4 <= __mul_41_stream_ivalid_3;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_5 <= __mul_41_stream_ivalid_4;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_6 <= __mul_41_stream_ivalid_5;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_7 <= __mul_41_stream_ivalid_6;
      end 
      if(_mul_41_stream_oready) begin
        __mul_41_stream_ivalid_8 <= __mul_41_stream_ivalid_7;
      end 
      if(_mul_41_stream_oready) begin
        _greaterthan_data_872 <= mul_41_rshift_data > 1'sd0;
      end 
      if(_mul_41_stream_oready) begin
        _minus_data_874 <= mul_41_rshift_data - 2'sd1;
      end 
      if(_mul_41_stream_oready) begin
        _greatereq_data_885 <= mul_41_x_data >= 1'sd0;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2323__variable_869 <= mul_41_x_data;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2326__variable_870 <= mul_41_y_data;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2329__variable_871 <= mul_41_rshift_data;
      end 
      if(_mul_41_stream_oready) begin
        _sll_data_876 <= 2'sd1 << _minus_data_874;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2320_greaterthan_872 <= _greaterthan_data_872;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2321_greatereq_885 <= _greatereq_data_885;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2324__delay_2323__variable_869 <= __delay_data_2323__variable_869;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2327__delay_2326__variable_870 <= __delay_data_2326__variable_870;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2330__delay_2329__variable_871 <= __delay_data_2329__variable_871;
      end 
      if(_mul_41_stream_oready) begin
        _cond_data_882 <= (__delay_data_2320_greaterthan_872)? _sll_data_876 : 1'sd0;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2322__delay_2321_greatereq_885 <= __delay_data_2321_greatereq_885;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2325__delay_2324__delay_2323__variable_869 <= __delay_data_2324__delay_2323__variable_869;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2328__delay_2327__delay_2326__variable_870 <= __delay_data_2327__delay_2326__variable_870;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2331__delay_2330__delay_2329__variable_871 <= __delay_data_2330__delay_2329__variable_871;
      end 
      if(_mul_41_stream_oready) begin
        __muladd_madd_odata_reg_888 <= __muladd_madd_odata_888;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2332__delay_2331__delay_2330____variable_871 <= __delay_data_2331__delay_2330__delay_2329__variable_871;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2333__delay_2332__delay_2331____variable_871 <= __delay_data_2332__delay_2331__delay_2330____variable_871;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2334__delay_2333__delay_2332____variable_871 <= __delay_data_2333__delay_2332__delay_2331____variable_871;
      end 
      if(_mul_41_stream_oready) begin
        __delay_data_2335__delay_2334__delay_2333____variable_871 <= __delay_data_2334__delay_2333__delay_2332____variable_871;
      end 
      if(_mul_41_stream_oready) begin
        _sra_data_889 <= __muladd_data_888 >>> __delay_data_2335__delay_2334__delay_2333____variable_871;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_869 <= _cond_data_2200;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_870 <= _cond_data_1557;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_871 <= __delay_data_2924__delay_2923_plus_2336;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1695 <= _mul_41_source_start;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1696 <= _tmp_1695;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1697 <= _tmp_1696;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1698 <= _mul_41_source_start;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1699 <= _tmp_1698;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1700 <= _tmp_1699;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1701 <= _tmp_1700;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1702 <= _tmp_1701;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1703 <= _tmp_1702;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1704 <= _tmp_1703;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1705 <= _tmp_1704;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1706 <= _tmp_1705;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1707 <= _tmp_1706;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1708 <= _mul_41_source_stop;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1709 <= _tmp_1708;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1710 <= _tmp_1709;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1711 <= _tmp_1710;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1712 <= _tmp_1711;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1713 <= _tmp_1712;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1714 <= _tmp_1713;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1715 <= _tmp_1714;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1716 <= _tmp_1715;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1717 <= _tmp_1716;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1718 <= _mul_41_source_busy;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1719 <= _tmp_1718;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1720 <= _tmp_1719;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1721 <= _tmp_1720;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1722 <= _tmp_1721;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1723 <= _tmp_1722;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1724 <= _tmp_1723;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1725 <= _tmp_1724;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1726 <= _tmp_1725;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1727 <= _tmp_1726;
      end 
      if(_mul_41_stream_oready) begin
        _tmp_1728 <= _mul_41_sink_busy;
      end 
      if(!_mul_41_sink_busy && _tmp_1728) begin
        _mul_41_busy_reg <= 0;
      end 
      if(_mul_41_source_busy) begin
        _mul_41_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_41_fsm_1 = 1;
  localparam _mul_41_fsm_2 = 2;
  localparam _mul_41_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_41_fsm <= _mul_41_fsm_init;
      _mul_41_source_start <= 0;
      _mul_41_source_busy <= 0;
      _mul_41_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_41_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_41_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_41_stream_oready && _tmp_1697) begin
        _mul_41_stream_ivalid <= 1;
      end 
      if(_mul_41_stream_oready && 1'd0) begin
        _mul_41_stream_ivalid <= 0;
      end 
      case(_mul_41_fsm)
        _mul_41_fsm_init: begin
          if(_mul_41_run_flag) begin
            _mul_41_source_start <= 1;
          end 
          if(_mul_41_run_flag) begin
            _mul_41_fsm <= _mul_41_fsm_1;
          end 
        end
        _mul_41_fsm_1: begin
          if(_mul_41_source_start && _mul_41_stream_oready) begin
            _mul_41_source_start <= 0;
            _mul_41_source_busy <= 1;
          end 
          if(_mul_41_source_start && _mul_41_stream_oready) begin
            _mul_41_fsm <= _mul_41_fsm_2;
          end 
        end
        _mul_41_fsm_2: begin
          if(_mul_41_stream_oready) begin
            _mul_41_fsm <= _mul_41_fsm_3;
          end 
        end
        _mul_41_fsm_3: begin
          if(_mul_41_stream_oready && 1'd0) begin
            _mul_41_source_busy <= 0;
          end 
          if(_mul_41_stream_oready && 1'd0 && _mul_41_run_flag) begin
            _mul_41_source_start <= 1;
          end 
          if(_mul_41_stream_oready && 1'd0) begin
            _mul_41_fsm <= _mul_41_fsm_init;
          end 
          if(_mul_41_stream_oready && 1'd0 && _mul_41_run_flag) begin
            _mul_41_fsm <= _mul_41_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_42_x_source_ram_renable <= 0;
      _mul_42_x_source_fifo_deq <= 0;
      _mul_42_x_idle <= 1;
      _mul_42_y_source_ram_renable <= 0;
      _mul_42_y_source_fifo_deq <= 0;
      _mul_42_y_idle <= 1;
      _mul_42_rshift_source_ram_renable <= 0;
      _mul_42_rshift_source_fifo_deq <= 0;
      _mul_42_rshift_idle <= 1;
      _mul_42_z_sink_wenable <= 0;
      _mul_42_z_sink_fifo_enq <= 0;
      __mul_42_stream_ivalid_1 <= 0;
      __mul_42_stream_ivalid_2 <= 0;
      __mul_42_stream_ivalid_3 <= 0;
      __mul_42_stream_ivalid_4 <= 0;
      __mul_42_stream_ivalid_5 <= 0;
      __mul_42_stream_ivalid_6 <= 0;
      __mul_42_stream_ivalid_7 <= 0;
      __mul_42_stream_ivalid_8 <= 0;
      _greaterthan_data_893 <= 0;
      _minus_data_895 <= 0;
      _greatereq_data_906 <= 0;
      __delay_data_2342__variable_890 <= 0;
      __delay_data_2345__variable_891 <= 0;
      __delay_data_2348__variable_892 <= 0;
      _sll_data_897 <= 0;
      __delay_data_2339_greaterthan_893 <= 0;
      __delay_data_2340_greatereq_906 <= 0;
      __delay_data_2343__delay_2342__variable_890 <= 0;
      __delay_data_2346__delay_2345__variable_891 <= 0;
      __delay_data_2349__delay_2348__variable_892 <= 0;
      _cond_data_903 <= 0;
      __delay_data_2341__delay_2340_greatereq_906 <= 0;
      __delay_data_2344__delay_2343__delay_2342__variable_890 <= 0;
      __delay_data_2347__delay_2346__delay_2345__variable_891 <= 0;
      __delay_data_2350__delay_2349__delay_2348__variable_892 <= 0;
      __muladd_madd_odata_reg_909 <= 0;
      __delay_data_2351__delay_2350__delay_2349____variable_892 <= 0;
      __delay_data_2352__delay_2351__delay_2350____variable_892 <= 0;
      __delay_data_2353__delay_2352__delay_2351____variable_892 <= 0;
      __delay_data_2354__delay_2353__delay_2352____variable_892 <= 0;
      _sra_data_910 <= 0;
      __variable_wdata_890 <= 0;
      __variable_wdata_891 <= 0;
      __variable_wdata_892 <= 0;
      _tmp_1729 <= 0;
      _tmp_1730 <= 0;
      _tmp_1731 <= 0;
      _tmp_1732 <= 0;
      _tmp_1733 <= 0;
      _tmp_1734 <= 0;
      _tmp_1735 <= 0;
      _tmp_1736 <= 0;
      _tmp_1737 <= 0;
      _tmp_1738 <= 0;
      _tmp_1739 <= 0;
      _tmp_1740 <= 0;
      _tmp_1741 <= 0;
      _tmp_1742 <= 0;
      _tmp_1743 <= 0;
      _tmp_1744 <= 0;
      _tmp_1745 <= 0;
      _tmp_1746 <= 0;
      _tmp_1747 <= 0;
      _tmp_1748 <= 0;
      _tmp_1749 <= 0;
      _tmp_1750 <= 0;
      _tmp_1751 <= 0;
      _tmp_1752 <= 0;
      _tmp_1753 <= 0;
      _tmp_1754 <= 0;
      _tmp_1755 <= 0;
      _tmp_1756 <= 0;
      _tmp_1757 <= 0;
      _tmp_1758 <= 0;
      _tmp_1759 <= 0;
      _tmp_1760 <= 0;
      _tmp_1761 <= 0;
      _tmp_1762 <= 0;
      _mul_42_busy_reg <= 0;
    end else begin
      if(_mul_42_stream_oready) begin
        _mul_42_x_source_ram_renable <= 0;
        _mul_42_x_source_fifo_deq <= 0;
      end 
      _mul_42_x_idle <= _mul_42_x_idle;
      if(_mul_42_stream_oready) begin
        _mul_42_y_source_ram_renable <= 0;
        _mul_42_y_source_fifo_deq <= 0;
      end 
      _mul_42_y_idle <= _mul_42_y_idle;
      if(_mul_42_stream_oready) begin
        _mul_42_rshift_source_ram_renable <= 0;
        _mul_42_rshift_source_fifo_deq <= 0;
      end 
      _mul_42_rshift_idle <= _mul_42_rshift_idle;
      if(_mul_42_stream_oready) begin
        _mul_42_z_sink_wenable <= 0;
        _mul_42_z_sink_fifo_enq <= 0;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_1 <= _mul_42_stream_ivalid;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_2 <= __mul_42_stream_ivalid_1;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_3 <= __mul_42_stream_ivalid_2;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_4 <= __mul_42_stream_ivalid_3;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_5 <= __mul_42_stream_ivalid_4;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_6 <= __mul_42_stream_ivalid_5;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_7 <= __mul_42_stream_ivalid_6;
      end 
      if(_mul_42_stream_oready) begin
        __mul_42_stream_ivalid_8 <= __mul_42_stream_ivalid_7;
      end 
      if(_mul_42_stream_oready) begin
        _greaterthan_data_893 <= mul_42_rshift_data > 1'sd0;
      end 
      if(_mul_42_stream_oready) begin
        _minus_data_895 <= mul_42_rshift_data - 2'sd1;
      end 
      if(_mul_42_stream_oready) begin
        _greatereq_data_906 <= mul_42_x_data >= 1'sd0;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2342__variable_890 <= mul_42_x_data;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2345__variable_891 <= mul_42_y_data;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2348__variable_892 <= mul_42_rshift_data;
      end 
      if(_mul_42_stream_oready) begin
        _sll_data_897 <= 2'sd1 << _minus_data_895;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2339_greaterthan_893 <= _greaterthan_data_893;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2340_greatereq_906 <= _greatereq_data_906;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2343__delay_2342__variable_890 <= __delay_data_2342__variable_890;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2346__delay_2345__variable_891 <= __delay_data_2345__variable_891;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2349__delay_2348__variable_892 <= __delay_data_2348__variable_892;
      end 
      if(_mul_42_stream_oready) begin
        _cond_data_903 <= (__delay_data_2339_greaterthan_893)? _sll_data_897 : 1'sd0;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2341__delay_2340_greatereq_906 <= __delay_data_2340_greatereq_906;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2344__delay_2343__delay_2342__variable_890 <= __delay_data_2343__delay_2342__variable_890;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2347__delay_2346__delay_2345__variable_891 <= __delay_data_2346__delay_2345__variable_891;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2350__delay_2349__delay_2348__variable_892 <= __delay_data_2349__delay_2348__variable_892;
      end 
      if(_mul_42_stream_oready) begin
        __muladd_madd_odata_reg_909 <= __muladd_madd_odata_909;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2351__delay_2350__delay_2349____variable_892 <= __delay_data_2350__delay_2349__delay_2348__variable_892;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2352__delay_2351__delay_2350____variable_892 <= __delay_data_2351__delay_2350__delay_2349____variable_892;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2353__delay_2352__delay_2351____variable_892 <= __delay_data_2352__delay_2351__delay_2350____variable_892;
      end 
      if(_mul_42_stream_oready) begin
        __delay_data_2354__delay_2353__delay_2352____variable_892 <= __delay_data_2353__delay_2352__delay_2351____variable_892;
      end 
      if(_mul_42_stream_oready) begin
        _sra_data_910 <= __muladd_data_909 >>> __delay_data_2354__delay_2353__delay_2352____variable_892;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_890 <= _cond_data_2202;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_891 <= _cond_data_1559;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_892 <= __delay_data_2934__delay_2933_plus_2355;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1729 <= _mul_42_source_start;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1730 <= _tmp_1729;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1731 <= _tmp_1730;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1732 <= _mul_42_source_start;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1733 <= _tmp_1732;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1734 <= _tmp_1733;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1735 <= _tmp_1734;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1736 <= _tmp_1735;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1737 <= _tmp_1736;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1738 <= _tmp_1737;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1739 <= _tmp_1738;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1740 <= _tmp_1739;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1741 <= _tmp_1740;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1742 <= _mul_42_source_stop;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1743 <= _tmp_1742;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1744 <= _tmp_1743;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1745 <= _tmp_1744;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1746 <= _tmp_1745;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1747 <= _tmp_1746;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1748 <= _tmp_1747;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1749 <= _tmp_1748;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1750 <= _tmp_1749;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1751 <= _tmp_1750;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1752 <= _mul_42_source_busy;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1753 <= _tmp_1752;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1754 <= _tmp_1753;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1755 <= _tmp_1754;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1756 <= _tmp_1755;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1757 <= _tmp_1756;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1758 <= _tmp_1757;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1759 <= _tmp_1758;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1760 <= _tmp_1759;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1761 <= _tmp_1760;
      end 
      if(_mul_42_stream_oready) begin
        _tmp_1762 <= _mul_42_sink_busy;
      end 
      if(!_mul_42_sink_busy && _tmp_1762) begin
        _mul_42_busy_reg <= 0;
      end 
      if(_mul_42_source_busy) begin
        _mul_42_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_42_fsm_1 = 1;
  localparam _mul_42_fsm_2 = 2;
  localparam _mul_42_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_42_fsm <= _mul_42_fsm_init;
      _mul_42_source_start <= 0;
      _mul_42_source_busy <= 0;
      _mul_42_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_42_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_42_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_42_stream_oready && _tmp_1731) begin
        _mul_42_stream_ivalid <= 1;
      end 
      if(_mul_42_stream_oready && 1'd0) begin
        _mul_42_stream_ivalid <= 0;
      end 
      case(_mul_42_fsm)
        _mul_42_fsm_init: begin
          if(_mul_42_run_flag) begin
            _mul_42_source_start <= 1;
          end 
          if(_mul_42_run_flag) begin
            _mul_42_fsm <= _mul_42_fsm_1;
          end 
        end
        _mul_42_fsm_1: begin
          if(_mul_42_source_start && _mul_42_stream_oready) begin
            _mul_42_source_start <= 0;
            _mul_42_source_busy <= 1;
          end 
          if(_mul_42_source_start && _mul_42_stream_oready) begin
            _mul_42_fsm <= _mul_42_fsm_2;
          end 
        end
        _mul_42_fsm_2: begin
          if(_mul_42_stream_oready) begin
            _mul_42_fsm <= _mul_42_fsm_3;
          end 
        end
        _mul_42_fsm_3: begin
          if(_mul_42_stream_oready && 1'd0) begin
            _mul_42_source_busy <= 0;
          end 
          if(_mul_42_stream_oready && 1'd0 && _mul_42_run_flag) begin
            _mul_42_source_start <= 1;
          end 
          if(_mul_42_stream_oready && 1'd0) begin
            _mul_42_fsm <= _mul_42_fsm_init;
          end 
          if(_mul_42_stream_oready && 1'd0 && _mul_42_run_flag) begin
            _mul_42_fsm <= _mul_42_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_43_x_source_ram_renable <= 0;
      _mul_43_x_source_fifo_deq <= 0;
      _mul_43_x_idle <= 1;
      _mul_43_y_source_ram_renable <= 0;
      _mul_43_y_source_fifo_deq <= 0;
      _mul_43_y_idle <= 1;
      _mul_43_rshift_source_ram_renable <= 0;
      _mul_43_rshift_source_fifo_deq <= 0;
      _mul_43_rshift_idle <= 1;
      _mul_43_z_sink_wenable <= 0;
      _mul_43_z_sink_fifo_enq <= 0;
      __mul_43_stream_ivalid_1 <= 0;
      __mul_43_stream_ivalid_2 <= 0;
      __mul_43_stream_ivalid_3 <= 0;
      __mul_43_stream_ivalid_4 <= 0;
      __mul_43_stream_ivalid_5 <= 0;
      __mul_43_stream_ivalid_6 <= 0;
      __mul_43_stream_ivalid_7 <= 0;
      __mul_43_stream_ivalid_8 <= 0;
      _greaterthan_data_914 <= 0;
      _minus_data_916 <= 0;
      _greatereq_data_927 <= 0;
      __delay_data_2361__variable_911 <= 0;
      __delay_data_2364__variable_912 <= 0;
      __delay_data_2367__variable_913 <= 0;
      _sll_data_918 <= 0;
      __delay_data_2358_greaterthan_914 <= 0;
      __delay_data_2359_greatereq_927 <= 0;
      __delay_data_2362__delay_2361__variable_911 <= 0;
      __delay_data_2365__delay_2364__variable_912 <= 0;
      __delay_data_2368__delay_2367__variable_913 <= 0;
      _cond_data_924 <= 0;
      __delay_data_2360__delay_2359_greatereq_927 <= 0;
      __delay_data_2363__delay_2362__delay_2361__variable_911 <= 0;
      __delay_data_2366__delay_2365__delay_2364__variable_912 <= 0;
      __delay_data_2369__delay_2368__delay_2367__variable_913 <= 0;
      __muladd_madd_odata_reg_930 <= 0;
      __delay_data_2370__delay_2369__delay_2368____variable_913 <= 0;
      __delay_data_2371__delay_2370__delay_2369____variable_913 <= 0;
      __delay_data_2372__delay_2371__delay_2370____variable_913 <= 0;
      __delay_data_2373__delay_2372__delay_2371____variable_913 <= 0;
      _sra_data_931 <= 0;
      __variable_wdata_911 <= 0;
      __variable_wdata_912 <= 0;
      __variable_wdata_913 <= 0;
      _tmp_1763 <= 0;
      _tmp_1764 <= 0;
      _tmp_1765 <= 0;
      _tmp_1766 <= 0;
      _tmp_1767 <= 0;
      _tmp_1768 <= 0;
      _tmp_1769 <= 0;
      _tmp_1770 <= 0;
      _tmp_1771 <= 0;
      _tmp_1772 <= 0;
      _tmp_1773 <= 0;
      _tmp_1774 <= 0;
      _tmp_1775 <= 0;
      _tmp_1776 <= 0;
      _tmp_1777 <= 0;
      _tmp_1778 <= 0;
      _tmp_1779 <= 0;
      _tmp_1780 <= 0;
      _tmp_1781 <= 0;
      _tmp_1782 <= 0;
      _tmp_1783 <= 0;
      _tmp_1784 <= 0;
      _tmp_1785 <= 0;
      _tmp_1786 <= 0;
      _tmp_1787 <= 0;
      _tmp_1788 <= 0;
      _tmp_1789 <= 0;
      _tmp_1790 <= 0;
      _tmp_1791 <= 0;
      _tmp_1792 <= 0;
      _tmp_1793 <= 0;
      _tmp_1794 <= 0;
      _tmp_1795 <= 0;
      _tmp_1796 <= 0;
      _mul_43_busy_reg <= 0;
    end else begin
      if(_mul_43_stream_oready) begin
        _mul_43_x_source_ram_renable <= 0;
        _mul_43_x_source_fifo_deq <= 0;
      end 
      _mul_43_x_idle <= _mul_43_x_idle;
      if(_mul_43_stream_oready) begin
        _mul_43_y_source_ram_renable <= 0;
        _mul_43_y_source_fifo_deq <= 0;
      end 
      _mul_43_y_idle <= _mul_43_y_idle;
      if(_mul_43_stream_oready) begin
        _mul_43_rshift_source_ram_renable <= 0;
        _mul_43_rshift_source_fifo_deq <= 0;
      end 
      _mul_43_rshift_idle <= _mul_43_rshift_idle;
      if(_mul_43_stream_oready) begin
        _mul_43_z_sink_wenable <= 0;
        _mul_43_z_sink_fifo_enq <= 0;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_1 <= _mul_43_stream_ivalid;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_2 <= __mul_43_stream_ivalid_1;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_3 <= __mul_43_stream_ivalid_2;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_4 <= __mul_43_stream_ivalid_3;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_5 <= __mul_43_stream_ivalid_4;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_6 <= __mul_43_stream_ivalid_5;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_7 <= __mul_43_stream_ivalid_6;
      end 
      if(_mul_43_stream_oready) begin
        __mul_43_stream_ivalid_8 <= __mul_43_stream_ivalid_7;
      end 
      if(_mul_43_stream_oready) begin
        _greaterthan_data_914 <= mul_43_rshift_data > 1'sd0;
      end 
      if(_mul_43_stream_oready) begin
        _minus_data_916 <= mul_43_rshift_data - 2'sd1;
      end 
      if(_mul_43_stream_oready) begin
        _greatereq_data_927 <= mul_43_x_data >= 1'sd0;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2361__variable_911 <= mul_43_x_data;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2364__variable_912 <= mul_43_y_data;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2367__variable_913 <= mul_43_rshift_data;
      end 
      if(_mul_43_stream_oready) begin
        _sll_data_918 <= 2'sd1 << _minus_data_916;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2358_greaterthan_914 <= _greaterthan_data_914;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2359_greatereq_927 <= _greatereq_data_927;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2362__delay_2361__variable_911 <= __delay_data_2361__variable_911;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2365__delay_2364__variable_912 <= __delay_data_2364__variable_912;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2368__delay_2367__variable_913 <= __delay_data_2367__variable_913;
      end 
      if(_mul_43_stream_oready) begin
        _cond_data_924 <= (__delay_data_2358_greaterthan_914)? _sll_data_918 : 1'sd0;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2360__delay_2359_greatereq_927 <= __delay_data_2359_greatereq_927;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2363__delay_2362__delay_2361__variable_911 <= __delay_data_2362__delay_2361__variable_911;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2366__delay_2365__delay_2364__variable_912 <= __delay_data_2365__delay_2364__variable_912;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2369__delay_2368__delay_2367__variable_913 <= __delay_data_2368__delay_2367__variable_913;
      end 
      if(_mul_43_stream_oready) begin
        __muladd_madd_odata_reg_930 <= __muladd_madd_odata_930;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2370__delay_2369__delay_2368____variable_913 <= __delay_data_2369__delay_2368__delay_2367__variable_913;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2371__delay_2370__delay_2369____variable_913 <= __delay_data_2370__delay_2369__delay_2368____variable_913;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2372__delay_2371__delay_2370____variable_913 <= __delay_data_2371__delay_2370__delay_2369____variable_913;
      end 
      if(_mul_43_stream_oready) begin
        __delay_data_2373__delay_2372__delay_2371____variable_913 <= __delay_data_2372__delay_2371__delay_2370____variable_913;
      end 
      if(_mul_43_stream_oready) begin
        _sra_data_931 <= __muladd_data_930 >>> __delay_data_2373__delay_2372__delay_2371____variable_913;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_911 <= _cond_data_2204;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_912 <= _cond_data_1561;
      end 
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_913 <= __delay_data_2944__delay_2943_plus_2374;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1763 <= _mul_43_source_start;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1764 <= _tmp_1763;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1765 <= _tmp_1764;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1766 <= _mul_43_source_start;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1767 <= _tmp_1766;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1768 <= _tmp_1767;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1769 <= _tmp_1768;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1770 <= _tmp_1769;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1771 <= _tmp_1770;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1772 <= _tmp_1771;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1773 <= _tmp_1772;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1774 <= _tmp_1773;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1775 <= _tmp_1774;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1776 <= _mul_43_source_stop;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1777 <= _tmp_1776;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1778 <= _tmp_1777;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1779 <= _tmp_1778;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1780 <= _tmp_1779;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1781 <= _tmp_1780;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1782 <= _tmp_1781;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1783 <= _tmp_1782;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1784 <= _tmp_1783;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1785 <= _tmp_1784;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1786 <= _mul_43_source_busy;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1787 <= _tmp_1786;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1788 <= _tmp_1787;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1789 <= _tmp_1788;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1790 <= _tmp_1789;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1791 <= _tmp_1790;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1792 <= _tmp_1791;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1793 <= _tmp_1792;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1794 <= _tmp_1793;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1795 <= _tmp_1794;
      end 
      if(_mul_43_stream_oready) begin
        _tmp_1796 <= _mul_43_sink_busy;
      end 
      if(!_mul_43_sink_busy && _tmp_1796) begin
        _mul_43_busy_reg <= 0;
      end 
      if(_mul_43_source_busy) begin
        _mul_43_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_43_fsm_1 = 1;
  localparam _mul_43_fsm_2 = 2;
  localparam _mul_43_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_43_fsm <= _mul_43_fsm_init;
      _mul_43_source_start <= 0;
      _mul_43_source_busy <= 0;
      _mul_43_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_3 && _stream_conv2d_4_stream_oready) begin
        _mul_43_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_43_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_43_stream_oready && _tmp_1765) begin
        _mul_43_stream_ivalid <= 1;
      end 
      if(_mul_43_stream_oready && 1'd0) begin
        _mul_43_stream_ivalid <= 0;
      end 
      case(_mul_43_fsm)
        _mul_43_fsm_init: begin
          if(_mul_43_run_flag) begin
            _mul_43_source_start <= 1;
          end 
          if(_mul_43_run_flag) begin
            _mul_43_fsm <= _mul_43_fsm_1;
          end 
        end
        _mul_43_fsm_1: begin
          if(_mul_43_source_start && _mul_43_stream_oready) begin
            _mul_43_source_start <= 0;
            _mul_43_source_busy <= 1;
          end 
          if(_mul_43_source_start && _mul_43_stream_oready) begin
            _mul_43_fsm <= _mul_43_fsm_2;
          end 
        end
        _mul_43_fsm_2: begin
          if(_mul_43_stream_oready) begin
            _mul_43_fsm <= _mul_43_fsm_3;
          end 
        end
        _mul_43_fsm_3: begin
          if(_mul_43_stream_oready && 1'd0) begin
            _mul_43_source_busy <= 0;
          end 
          if(_mul_43_stream_oready && 1'd0 && _mul_43_run_flag) begin
            _mul_43_source_start <= 1;
          end 
          if(_mul_43_stream_oready && 1'd0) begin
            _mul_43_fsm <= _mul_43_fsm_init;
          end 
          if(_mul_43_stream_oready && 1'd0 && _mul_43_run_flag) begin
            _mul_43_fsm <= _mul_43_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_44_x_source_ram_renable <= 0;
      __reduce_max_44_x_source_fifo_deq <= 0;
      __reduce_max_44_x_idle <= 1;
      __reduce_max_44_data_sink_wenable <= 0;
      __reduce_max_44_data_sink_fifo_enq <= 0;
      __reduce_max_44_valid_sink_wenable <= 0;
      __reduce_max_44_valid_sink_fifo_enq <= 0;
      ___reduce_max_44_stream_ivalid_1 <= 0;
      _reducemax_data_935 <= -17'sd32768;
      _reducemax_count_935 <= 0;
      _reducemax_prev_count_max_935 <= 0;
      _pulse_data_937 <= 1'sd0;
      _pulse_count_937 <= 0;
      _pulse_prev_count_max_937 <= 0;
      __variable_wdata_934 <= 0;
      __variable_wdata_932 <= 0;
      __variable_wdata_933 <= 0;
      _tmp_2083 <= 0;
      _tmp_2084 <= 0;
      _tmp_2085 <= 0;
      _tmp_2086 <= 0;
      _tmp_2087 <= 0;
      _tmp_2088 <= 0;
      _tmp_2089 <= 0;
      _tmp_2090 <= 0;
      _tmp_2091 <= 0;
      _tmp_2092 <= 0;
      _tmp_2093 <= 0;
      _tmp_2094 <= 0;
      _tmp_2095 <= 0;
      _tmp_2096 <= 0;
      _tmp_2097 <= 0;
      _tmp_2098 <= 0;
      _tmp_2099 <= 0;
      _tmp_2100 <= 0;
      _tmp_2101 <= 0;
      _tmp_2102 <= 0;
      __reduce_max_44_busy_reg <= 0;
    end else begin
      if(__reduce_max_44_stream_oready) begin
        __reduce_max_44_x_source_ram_renable <= 0;
        __reduce_max_44_x_source_fifo_deq <= 0;
      end 
      __reduce_max_44_x_idle <= __reduce_max_44_x_idle;
      if(__reduce_max_44_stream_oready) begin
        __reduce_max_44_data_sink_wenable <= 0;
        __reduce_max_44_data_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_44_stream_oready) begin
        __reduce_max_44_valid_sink_wenable <= 0;
        __reduce_max_44_valid_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_44_stream_oready) begin
        ___reduce_max_44_stream_ivalid_1 <= __reduce_max_44_stream_ivalid;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready && _reducemax_reset_cond_935) begin
        _reducemax_data_935 <= -17'sd32768;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready) begin
        _reducemax_count_935 <= (_reducemax_current_count_935 >= _reduce_max_44_size_data - 1)? 0 : _reducemax_current_count_935 + 1;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready) begin
        _reducemax_prev_count_max_935 <= _reducemax_current_count_935 >= _reduce_max_44_size_data - 1;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready) begin
        _reducemax_data_935 <= (_reducemax_current_data_935 < _reduce_max_44_x_data)? _reduce_max_44_x_data : _reducemax_current_data_935;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready && _pulse_reset_cond_937) begin
        _pulse_data_937 <= 1'sd0;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready) begin
        _pulse_count_937 <= (_pulse_current_count_937 >= _reduce_max_44_size_data - 1)? 0 : _pulse_current_count_937 + 1;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready) begin
        _pulse_prev_count_max_937 <= _pulse_current_count_937 >= _reduce_max_44_size_data - 1;
      end 
      if(__reduce_max_44_stream_ivalid && __reduce_max_44_stream_oready) begin
        _pulse_data_937 <= _pulse_current_count_937 >= _reduce_max_44_size_data - 1;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_934 <= __delay_data_3113__delay_3112__delay_3111__variable_2420;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_932 <= _cond_data_2434;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_933 <= __delay_data_3116__delay_3115__delay_3114__variable_2417;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2083 <= __reduce_max_44_source_start;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2084 <= _tmp_2083;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2085 <= _tmp_2084;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2086 <= __reduce_max_44_source_start;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2087 <= _tmp_2086;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2088 <= _tmp_2087;
      end 
      if(__reduce_max_44_stream_oready && _tmp_2088) begin
        __variable_wdata_934 <= 1;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2089 <= __reduce_max_44_source_start;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2090 <= _tmp_2089;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2091 <= _tmp_2090;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2092 <= _tmp_2091;
      end 
      if(__reduce_max_44_stream_oready && _tmp_2092) begin
        __variable_wdata_934 <= 0;
      end 
      if(__reduce_max_44_stream_oready && 1'd0) begin
        __variable_wdata_934 <= 1;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2093 <= __reduce_max_44_source_start;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2094 <= _tmp_2093;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2095 <= _tmp_2094;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2096 <= __reduce_max_44_source_stop;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2097 <= _tmp_2096;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2098 <= _tmp_2097;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2099 <= __reduce_max_44_source_busy;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2100 <= _tmp_2099;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2101 <= _tmp_2100;
      end 
      if(__reduce_max_44_stream_oready) begin
        _tmp_2102 <= __reduce_max_44_sink_busy;
      end 
      if(!__reduce_max_44_sink_busy && _tmp_2102) begin
        __reduce_max_44_busy_reg <= 0;
      end 
      if(__reduce_max_44_source_busy) begin
        __reduce_max_44_busy_reg <= 1;
      end 
    end
  end

  localparam __reduce_max_44_fsm_1 = 1;
  localparam __reduce_max_44_fsm_2 = 2;
  localparam __reduce_max_44_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_44_fsm <= __reduce_max_44_fsm_init;
      __reduce_max_44_source_start <= 0;
      __reduce_max_44_source_busy <= 0;
      __reduce_max_44_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __reduce_max_44_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_busy) begin
        __reduce_max_44_source_busy <= _stream_max_pool_serial_6_source_busy;
      end 
      if(__reduce_max_44_stream_oready && _tmp_2085) begin
        __reduce_max_44_stream_ivalid <= 1;
      end 
      if(__reduce_max_44_stream_oready && 1'd0) begin
        __reduce_max_44_stream_ivalid <= 0;
      end 
      case(__reduce_max_44_fsm)
        __reduce_max_44_fsm_init: begin
          if(__reduce_max_44_run_flag) begin
            __reduce_max_44_source_start <= 1;
          end 
          if(__reduce_max_44_run_flag) begin
            __reduce_max_44_fsm <= __reduce_max_44_fsm_1;
          end 
        end
        __reduce_max_44_fsm_1: begin
          if(__reduce_max_44_source_start && __reduce_max_44_stream_oready) begin
            __reduce_max_44_source_start <= 0;
            __reduce_max_44_source_busy <= 1;
          end 
          if(__reduce_max_44_source_start && __reduce_max_44_stream_oready) begin
            __reduce_max_44_fsm <= __reduce_max_44_fsm_2;
          end 
        end
        __reduce_max_44_fsm_2: begin
          if(__reduce_max_44_stream_oready) begin
            __reduce_max_44_fsm <= __reduce_max_44_fsm_3;
          end 
        end
        __reduce_max_44_fsm_3: begin
          if(__reduce_max_44_stream_oready && 1'd0) begin
            __reduce_max_44_source_busy <= 0;
          end 
          if(__reduce_max_44_stream_oready && 1'd0 && __reduce_max_44_run_flag) begin
            __reduce_max_44_source_start <= 1;
          end 
          if(__reduce_max_44_stream_oready && 1'd0) begin
            __reduce_max_44_fsm <= __reduce_max_44_fsm_init;
          end 
          if(__reduce_max_44_stream_oready && 1'd0 && __reduce_max_44_run_flag) begin
            __reduce_max_44_fsm <= __reduce_max_44_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_45_x_source_ram_renable <= 0;
      __reduce_max_45_x_source_fifo_deq <= 0;
      __reduce_max_45_x_idle <= 1;
      __reduce_max_45_data_sink_wenable <= 0;
      __reduce_max_45_data_sink_fifo_enq <= 0;
      __reduce_max_45_valid_sink_wenable <= 0;
      __reduce_max_45_valid_sink_fifo_enq <= 0;
      ___reduce_max_45_stream_ivalid_1 <= 0;
      _reducemax_data_942 <= -17'sd32768;
      _reducemax_count_942 <= 0;
      _reducemax_prev_count_max_942 <= 0;
      _pulse_data_944 <= 1'sd0;
      _pulse_count_944 <= 0;
      _pulse_prev_count_max_944 <= 0;
      __variable_wdata_941 <= 0;
      __variable_wdata_939 <= 0;
      __variable_wdata_940 <= 0;
      _tmp_2103 <= 0;
      _tmp_2104 <= 0;
      _tmp_2105 <= 0;
      _tmp_2106 <= 0;
      _tmp_2107 <= 0;
      _tmp_2108 <= 0;
      _tmp_2109 <= 0;
      _tmp_2110 <= 0;
      _tmp_2111 <= 0;
      _tmp_2112 <= 0;
      _tmp_2113 <= 0;
      _tmp_2114 <= 0;
      _tmp_2115 <= 0;
      _tmp_2116 <= 0;
      _tmp_2117 <= 0;
      _tmp_2118 <= 0;
      _tmp_2119 <= 0;
      _tmp_2120 <= 0;
      _tmp_2121 <= 0;
      _tmp_2122 <= 0;
      __reduce_max_45_busy_reg <= 0;
    end else begin
      if(__reduce_max_45_stream_oready) begin
        __reduce_max_45_x_source_ram_renable <= 0;
        __reduce_max_45_x_source_fifo_deq <= 0;
      end 
      __reduce_max_45_x_idle <= __reduce_max_45_x_idle;
      if(__reduce_max_45_stream_oready) begin
        __reduce_max_45_data_sink_wenable <= 0;
        __reduce_max_45_data_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_45_stream_oready) begin
        __reduce_max_45_valid_sink_wenable <= 0;
        __reduce_max_45_valid_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_45_stream_oready) begin
        ___reduce_max_45_stream_ivalid_1 <= __reduce_max_45_stream_ivalid;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready && _reducemax_reset_cond_942) begin
        _reducemax_data_942 <= -17'sd32768;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready) begin
        _reducemax_count_942 <= (_reducemax_current_count_942 >= _reduce_max_45_size_data - 1)? 0 : _reducemax_current_count_942 + 1;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready) begin
        _reducemax_prev_count_max_942 <= _reducemax_current_count_942 >= _reduce_max_45_size_data - 1;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready) begin
        _reducemax_data_942 <= (_reducemax_current_data_942 < _reduce_max_45_x_data)? _reduce_max_45_x_data : _reducemax_current_data_942;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready && _pulse_reset_cond_944) begin
        _pulse_data_944 <= 1'sd0;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready) begin
        _pulse_count_944 <= (_pulse_current_count_944 >= _reduce_max_45_size_data - 1)? 0 : _pulse_current_count_944 + 1;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready) begin
        _pulse_prev_count_max_944 <= _pulse_current_count_944 >= _reduce_max_45_size_data - 1;
      end 
      if(__reduce_max_45_stream_ivalid && __reduce_max_45_stream_oready) begin
        _pulse_data_944 <= _pulse_current_count_944 >= _reduce_max_45_size_data - 1;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_941 <= __delay_data_3113__delay_3112__delay_3111__variable_2420;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_939 <= _cond_data_2439;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_940 <= __delay_data_3116__delay_3115__delay_3114__variable_2417;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2103 <= __reduce_max_45_source_start;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2104 <= _tmp_2103;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2105 <= _tmp_2104;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2106 <= __reduce_max_45_source_start;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2107 <= _tmp_2106;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2108 <= _tmp_2107;
      end 
      if(__reduce_max_45_stream_oready && _tmp_2108) begin
        __variable_wdata_941 <= 1;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2109 <= __reduce_max_45_source_start;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2110 <= _tmp_2109;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2111 <= _tmp_2110;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2112 <= _tmp_2111;
      end 
      if(__reduce_max_45_stream_oready && _tmp_2112) begin
        __variable_wdata_941 <= 0;
      end 
      if(__reduce_max_45_stream_oready && 1'd0) begin
        __variable_wdata_941 <= 1;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2113 <= __reduce_max_45_source_start;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2114 <= _tmp_2113;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2115 <= _tmp_2114;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2116 <= __reduce_max_45_source_stop;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2117 <= _tmp_2116;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2118 <= _tmp_2117;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2119 <= __reduce_max_45_source_busy;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2120 <= _tmp_2119;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2121 <= _tmp_2120;
      end 
      if(__reduce_max_45_stream_oready) begin
        _tmp_2122 <= __reduce_max_45_sink_busy;
      end 
      if(!__reduce_max_45_sink_busy && _tmp_2122) begin
        __reduce_max_45_busy_reg <= 0;
      end 
      if(__reduce_max_45_source_busy) begin
        __reduce_max_45_busy_reg <= 1;
      end 
    end
  end

  localparam __reduce_max_45_fsm_1 = 1;
  localparam __reduce_max_45_fsm_2 = 2;
  localparam __reduce_max_45_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_45_fsm <= __reduce_max_45_fsm_init;
      __reduce_max_45_source_start <= 0;
      __reduce_max_45_source_busy <= 0;
      __reduce_max_45_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __reduce_max_45_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_busy) begin
        __reduce_max_45_source_busy <= _stream_max_pool_serial_6_source_busy;
      end 
      if(__reduce_max_45_stream_oready && _tmp_2105) begin
        __reduce_max_45_stream_ivalid <= 1;
      end 
      if(__reduce_max_45_stream_oready && 1'd0) begin
        __reduce_max_45_stream_ivalid <= 0;
      end 
      case(__reduce_max_45_fsm)
        __reduce_max_45_fsm_init: begin
          if(__reduce_max_45_run_flag) begin
            __reduce_max_45_source_start <= 1;
          end 
          if(__reduce_max_45_run_flag) begin
            __reduce_max_45_fsm <= __reduce_max_45_fsm_1;
          end 
        end
        __reduce_max_45_fsm_1: begin
          if(__reduce_max_45_source_start && __reduce_max_45_stream_oready) begin
            __reduce_max_45_source_start <= 0;
            __reduce_max_45_source_busy <= 1;
          end 
          if(__reduce_max_45_source_start && __reduce_max_45_stream_oready) begin
            __reduce_max_45_fsm <= __reduce_max_45_fsm_2;
          end 
        end
        __reduce_max_45_fsm_2: begin
          if(__reduce_max_45_stream_oready) begin
            __reduce_max_45_fsm <= __reduce_max_45_fsm_3;
          end 
        end
        __reduce_max_45_fsm_3: begin
          if(__reduce_max_45_stream_oready && 1'd0) begin
            __reduce_max_45_source_busy <= 0;
          end 
          if(__reduce_max_45_stream_oready && 1'd0 && __reduce_max_45_run_flag) begin
            __reduce_max_45_source_start <= 1;
          end 
          if(__reduce_max_45_stream_oready && 1'd0) begin
            __reduce_max_45_fsm <= __reduce_max_45_fsm_init;
          end 
          if(__reduce_max_45_stream_oready && 1'd0 && __reduce_max_45_run_flag) begin
            __reduce_max_45_fsm <= __reduce_max_45_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_7_source_ram_renable <= 0;
      _stream_conv2d_4_source_7_source_fifo_deq <= 0;
      _stream_conv2d_4_source_7_idle <= 1;
      _stream_conv2d_4_source_9_source_ram_renable <= 0;
      _stream_conv2d_4_source_9_source_fifo_deq <= 0;
      _stream_conv2d_4_source_9_idle <= 1;
      _stream_conv2d_4_source_11_source_ram_renable <= 0;
      _stream_conv2d_4_source_11_source_fifo_deq <= 0;
      _stream_conv2d_4_source_11_idle <= 1;
      _stream_conv2d_4_source_13_source_ram_renable <= 0;
      _stream_conv2d_4_source_13_source_fifo_deq <= 0;
      _stream_conv2d_4_source_13_idle <= 1;
      _stream_conv2d_4_source_15_source_ram_renable <= 0;
      _stream_conv2d_4_source_15_source_fifo_deq <= 0;
      _stream_conv2d_4_source_15_idle <= 1;
      _stream_conv2d_4_source_20_source_ram_renable <= 0;
      _stream_conv2d_4_source_20_source_fifo_deq <= 0;
      _stream_conv2d_4_source_20_idle <= 1;
      _stream_conv2d_4_source_21_source_ram_renable <= 0;
      _stream_conv2d_4_source_21_source_fifo_deq <= 0;
      _stream_conv2d_4_source_21_idle <= 1;
      _stream_conv2d_4_source_22_source_ram_renable <= 0;
      _stream_conv2d_4_source_22_source_fifo_deq <= 0;
      _stream_conv2d_4_source_22_idle <= 1;
      _stream_conv2d_4_source_23_source_ram_renable <= 0;
      _stream_conv2d_4_source_23_source_fifo_deq <= 0;
      _stream_conv2d_4_source_23_idle <= 1;
      _stream_conv2d_4_source_24_source_ram_renable <= 0;
      _stream_conv2d_4_source_24_source_fifo_deq <= 0;
      _stream_conv2d_4_source_24_idle <= 1;
      _stream_conv2d_4_source_25_source_ram_renable <= 0;
      _stream_conv2d_4_source_25_source_fifo_deq <= 0;
      _stream_conv2d_4_source_25_idle <= 1;
      _stream_conv2d_4_source_26_source_ram_renable <= 0;
      _stream_conv2d_4_source_26_source_fifo_deq <= 0;
      _stream_conv2d_4_source_26_idle <= 1;
      _stream_conv2d_4_source_27_source_ram_renable <= 0;
      _stream_conv2d_4_source_27_source_fifo_deq <= 0;
      _stream_conv2d_4_source_27_idle <= 1;
      _stream_conv2d_4_source_28_source_ram_renable <= 0;
      _stream_conv2d_4_source_28_source_fifo_deq <= 0;
      _stream_conv2d_4_source_28_idle <= 1;
      _stream_conv2d_4_source_29_source_ram_renable <= 0;
      _stream_conv2d_4_source_29_source_fifo_deq <= 0;
      _stream_conv2d_4_source_29_idle <= 1;
      _stream_conv2d_4_source_30_source_ram_renable <= 0;
      _stream_conv2d_4_source_30_source_fifo_deq <= 0;
      _stream_conv2d_4_source_30_idle <= 1;
      _stream_conv2d_4_source_31_source_ram_renable <= 0;
      _stream_conv2d_4_source_31_source_fifo_deq <= 0;
      _stream_conv2d_4_source_31_idle <= 1;
      _stream_conv2d_4_source_32_source_ram_renable <= 0;
      _stream_conv2d_4_source_32_source_fifo_deq <= 0;
      _stream_conv2d_4_source_32_idle <= 1;
      _stream_conv2d_4_source_33_source_ram_renable <= 0;
      _stream_conv2d_4_source_33_source_fifo_deq <= 0;
      _stream_conv2d_4_source_33_idle <= 1;
      _stream_conv2d_4_source_34_source_ram_renable <= 0;
      _stream_conv2d_4_source_34_source_fifo_deq <= 0;
      _stream_conv2d_4_source_34_idle <= 1;
      _stream_conv2d_4_source_35_source_ram_renable <= 0;
      _stream_conv2d_4_source_35_source_fifo_deq <= 0;
      _stream_conv2d_4_source_35_idle <= 1;
      _stream_conv2d_4_source_36_source_ram_renable <= 0;
      _stream_conv2d_4_source_36_source_fifo_deq <= 0;
      _stream_conv2d_4_source_36_idle <= 1;
      _stream_conv2d_4_source_37_source_ram_renable <= 0;
      _stream_conv2d_4_source_37_source_fifo_deq <= 0;
      _stream_conv2d_4_source_37_idle <= 1;
      _stream_conv2d_4_source_38_source_ram_renable <= 0;
      _stream_conv2d_4_source_38_source_fifo_deq <= 0;
      _stream_conv2d_4_source_38_idle <= 1;
      _stream_conv2d_4_source_39_source_ram_renable <= 0;
      _stream_conv2d_4_source_39_source_fifo_deq <= 0;
      _stream_conv2d_4_source_39_idle <= 1;
      _stream_conv2d_4_source_40_source_ram_renable <= 0;
      _stream_conv2d_4_source_40_source_fifo_deq <= 0;
      _stream_conv2d_4_source_40_idle <= 1;
      _stream_conv2d_4_source_41_source_ram_renable <= 0;
      _stream_conv2d_4_source_41_source_fifo_deq <= 0;
      _stream_conv2d_4_source_41_idle <= 1;
      _stream_conv2d_4_source_42_source_ram_renable <= 0;
      _stream_conv2d_4_source_42_source_fifo_deq <= 0;
      _stream_conv2d_4_source_42_idle <= 1;
      _stream_conv2d_4_source_43_source_ram_renable <= 0;
      _stream_conv2d_4_source_43_source_fifo_deq <= 0;
      _stream_conv2d_4_source_43_idle <= 1;
      _stream_conv2d_4_source_44_source_ram_renable <= 0;
      _stream_conv2d_4_source_44_source_fifo_deq <= 0;
      _stream_conv2d_4_source_44_idle <= 1;
      _stream_conv2d_4_source_45_source_ram_renable <= 0;
      _stream_conv2d_4_source_45_source_fifo_deq <= 0;
      _stream_conv2d_4_source_45_idle <= 1;
      _stream_conv2d_4_source_46_source_ram_renable <= 0;
      _stream_conv2d_4_source_46_source_fifo_deq <= 0;
      _stream_conv2d_4_source_46_idle <= 1;
      _stream_conv2d_4_sink_89_sink_wenable <= 0;
      _stream_conv2d_4_sink_89_sink_fifo_enq <= 0;
      _stream_conv2d_4_sink_90_sink_wenable <= 0;
      _stream_conv2d_4_sink_90_sink_fifo_enq <= 0;
      __stream_conv2d_4_stream_ivalid_1 <= 0;
      __stream_conv2d_4_stream_ivalid_2 <= 0;
      __stream_conv2d_4_stream_ivalid_3 <= 0;
      __stream_conv2d_4_stream_ivalid_4 <= 0;
      __stream_conv2d_4_stream_ivalid_5 <= 0;
      __stream_conv2d_4_stream_ivalid_6 <= 0;
      __stream_conv2d_4_stream_ivalid_7 <= 0;
      __stream_conv2d_4_stream_ivalid_8 <= 0;
      __stream_conv2d_4_stream_ivalid_9 <= 0;
      __stream_conv2d_4_stream_ivalid_10 <= 0;
      __stream_conv2d_4_stream_ivalid_11 <= 0;
      __stream_conv2d_4_stream_ivalid_12 <= 0;
      __stream_conv2d_4_stream_ivalid_13 <= 0;
      __stream_conv2d_4_stream_ivalid_14 <= 0;
      __stream_conv2d_4_stream_ivalid_15 <= 0;
      __stream_conv2d_4_stream_ivalid_16 <= 0;
      __stream_conv2d_4_stream_ivalid_17 <= 0;
      __stream_conv2d_4_stream_ivalid_18 <= 0;
      __stream_conv2d_4_stream_ivalid_19 <= 0;
      __stream_conv2d_4_stream_ivalid_20 <= 0;
      __stream_conv2d_4_stream_ivalid_21 <= 0;
      __stream_conv2d_4_stream_ivalid_22 <= 0;
      __stream_conv2d_4_stream_ivalid_23 <= 0;
      __stream_conv2d_4_stream_ivalid_24 <= 0;
      __stream_conv2d_4_stream_ivalid_25 <= 0;
      __stream_conv2d_4_stream_ivalid_26 <= 0;
      __stream_conv2d_4_stream_ivalid_27 <= 0;
      __stream_conv2d_4_stream_ivalid_28 <= 0;
      __stream_conv2d_4_stream_ivalid_29 <= 0;
      __stream_conv2d_4_stream_ivalid_30 <= 0;
      __stream_conv2d_4_stream_ivalid_31 <= 0;
      __stream_conv2d_4_stream_ivalid_32 <= 0;
      __stream_conv2d_4_stream_ivalid_33 <= 0;
      __stream_conv2d_4_stream_ivalid_34 <= 0;
      _counter_data_952 <= 1'sd0;
      _counter_count_952 <= 1'sd0;
      _minus_data_957 <= 0;
      _minus_data_963 <= 0;
      _eq_data_1040 <= 0;
      _eq_data_1044 <= 0;
      _eq_data_1047 <= 0;
      _eq_data_1050 <= 0;
      _eq_data_1054 <= 0;
      _eq_data_1057 <= 0;
      _eq_data_1060 <= 0;
      _eq_data_1064 <= 0;
      _eq_data_1067 <= 0;
      _eq_data_1070 <= 0;
      _eq_data_1074 <= 0;
      _eq_data_1077 <= 0;
      _eq_data_1080 <= 0;
      _eq_data_1084 <= 0;
      _eq_data_1087 <= 0;
      _eq_data_1090 <= 0;
      _eq_data_1094 <= 0;
      _eq_data_1097 <= 0;
      _eq_data_1100 <= 0;
      _eq_data_1104 <= 0;
      _eq_data_1107 <= 0;
      _eq_data_1110 <= 0;
      _eq_data_1114 <= 0;
      _eq_data_1117 <= 0;
      _eq_data_1120 <= 0;
      _eq_data_1124 <= 0;
      _eq_data_1127 <= 0;
      _eq_data_1130 <= 0;
      _eq_data_1134 <= 0;
      _eq_data_1137 <= 0;
      _eq_data_1140 <= 0;
      _eq_data_1144 <= 0;
      _eq_data_1147 <= 0;
      _eq_data_1150 <= 0;
      _eq_data_1154 <= 0;
      _eq_data_1157 <= 0;
      _eq_data_1160 <= 0;
      _eq_data_1164 <= 0;
      _eq_data_1167 <= 0;
      _eq_data_1170 <= 0;
      _eq_data_1174 <= 0;
      _eq_data_1177 <= 0;
      _eq_data_1180 <= 0;
      _eq_data_1184 <= 0;
      _eq_data_1187 <= 0;
      _eq_data_1190 <= 0;
      _eq_data_1194 <= 0;
      _eq_data_1197 <= 0;
      _eq_data_1200 <= 0;
      _eq_data_1204 <= 0;
      _eq_data_1207 <= 0;
      _eq_data_1210 <= 0;
      _eq_data_1214 <= 0;
      _eq_data_1217 <= 0;
      _plus_data_1615 <= 0;
      _plus_data_1634 <= 0;
      _plus_data_1653 <= 0;
      _plus_data_1672 <= 0;
      _plus_data_1691 <= 0;
      _plus_data_1710 <= 0;
      _plus_data_1729 <= 0;
      _plus_data_1748 <= 0;
      _plus_data_1767 <= 0;
      _plus_data_1804 <= 0;
      _plus_data_1823 <= 0;
      _plus_data_1842 <= 0;
      _plus_data_1861 <= 0;
      _plus_data_1880 <= 0;
      _plus_data_1899 <= 0;
      _plus_data_1918 <= 0;
      _plus_data_1937 <= 0;
      _plus_data_1956 <= 0;
      _plus_data_1972 <= 0;
      _plus_data_1991 <= 0;
      _plus_data_2033 <= 0;
      _plus_data_2052 <= 0;
      _plus_data_2071 <= 0;
      _plus_data_2090 <= 0;
      _plus_data_2109 <= 0;
      _plus_data_2128 <= 0;
      _plus_data_2147 <= 0;
      _plus_data_2166 <= 0;
      _plus_data_2185 <= 0;
      _plus_data_2222 <= 0;
      _plus_data_2241 <= 0;
      _plus_data_2260 <= 0;
      _plus_data_2279 <= 0;
      _plus_data_2298 <= 0;
      _plus_data_2317 <= 0;
      _plus_data_2336 <= 0;
      _plus_data_2355 <= 0;
      _plus_data_2374 <= 0;
      _plus_data_2390 <= 0;
      _plus_data_2409 <= 0;
      __delay_data_2642_pointer_955 <= 0;
      __delay_data_2644__variable_1033 <= 0;
      __delay_data_2645__variable_1032 <= 0;
      __delay_data_2646__variable_1031 <= 0;
      __delay_data_2647__variable_1036 <= 0;
      __delay_data_2648__variable_1035 <= 0;
      __delay_data_2649__variable_1034 <= 0;
      __delay_data_2650__variable_1039 <= 0;
      __delay_data_2651__variable_1038 <= 0;
      __delay_data_2652__variable_1037 <= 0;
      __delay_data_2655_pointer_1562 <= 0;
      __delay_data_2658_reinterpretcast_1349 <= 0;
      __delay_data_2663_pointer_961 <= 0;
      __delay_data_2667_reinterpretcast_1353 <= 0;
      __delay_data_2674_pointer_1564 <= 0;
      __delay_data_2677_reinterpretcast_1357 <= 0;
      __delay_data_2684_reinterpretcast_1361 <= 0;
      __delay_data_2691_pointer_1566 <= 0;
      __delay_data_2694_reinterpretcast_1365 <= 0;
      __delay_data_2701_reinterpretcast_1369 <= 0;
      __delay_data_2708_pointer_1568 <= 0;
      __delay_data_2711_reinterpretcast_1373 <= 0;
      __delay_data_2718_reinterpretcast_1377 <= 0;
      __delay_data_2725_pointer_1570 <= 0;
      __delay_data_2728_reinterpretcast_1381 <= 0;
      __delay_data_2735_reinterpretcast_1385 <= 0;
      __delay_data_2742_pointer_1572 <= 0;
      __delay_data_2745_reinterpretcast_1389 <= 0;
      __delay_data_2752_reinterpretcast_1393 <= 0;
      __delay_data_2759_pointer_1574 <= 0;
      __delay_data_2762_reinterpretcast_1397 <= 0;
      __delay_data_2769_reinterpretcast_1401 <= 0;
      __delay_data_2776_pointer_1576 <= 0;
      __delay_data_2779_reinterpretcast_1405 <= 0;
      __delay_data_2786_reinterpretcast_1409 <= 0;
      __delay_data_2793_pointer_1578 <= 0;
      __delay_data_2796_reinterpretcast_1413 <= 0;
      __delay_data_2803_reinterpretcast_1417 <= 0;
      __delay_data_2808__variable_951 <= 0;
      __delay_data_2839__variable_946 <= 0;
      __delay_data_2855_reinterpretcast_1457 <= 0;
      __delay_data_2860_reinterpretcast_1461 <= 0;
      __delay_data_2865_reinterpretcast_1465 <= 0;
      __delay_data_2870_reinterpretcast_1469 <= 0;
      __delay_data_2875_reinterpretcast_1473 <= 0;
      __delay_data_2880_reinterpretcast_1477 <= 0;
      __delay_data_2885_reinterpretcast_1481 <= 0;
      __delay_data_2890_reinterpretcast_1485 <= 0;
      __delay_data_2895_reinterpretcast_1489 <= 0;
      __delay_data_2900_reinterpretcast_1493 <= 0;
      __delay_data_2905_reinterpretcast_1497 <= 0;
      __delay_data_2910_reinterpretcast_1501 <= 0;
      __delay_data_2915_reinterpretcast_1505 <= 0;
      __delay_data_2920_reinterpretcast_1509 <= 0;
      __delay_data_2925_reinterpretcast_1513 <= 0;
      __delay_data_2930_reinterpretcast_1517 <= 0;
      __delay_data_2935_reinterpretcast_1521 <= 0;
      __delay_data_2940_reinterpretcast_1525 <= 0;
      __delay_data_2960_cond_978 <= 0;
      __delay_data_2982_cond_990 <= 0;
      __delay_data_3028_cond_977 <= 0;
      __delay_data_3050_cond_989 <= 0;
      _eq_data_959 <= 0;
      _eq_data_965 <= 0;
      __delay_data_2643__delay_2642_pointer_955 <= 0;
      __delay_data_2653_reinterpretcast_1223 <= 0;
      __delay_data_2656__delay_2655_pointer_1562 <= 0;
      __delay_data_2659__delay_2658_reinterpretcast_1349 <= 0;
      __delay_data_2661_plus_1615 <= 0;
      __delay_data_2664__delay_2663_pointer_961 <= 0;
      __delay_data_2665_reinterpretcast_1227 <= 0;
      __delay_data_2668__delay_2667_reinterpretcast_1353 <= 0;
      __delay_data_2670_plus_1804 <= 0;
      __delay_data_2672_reinterpretcast_1231 <= 0;
      __delay_data_2675__delay_2674_pointer_1564 <= 0;
      __delay_data_2678__delay_2677_reinterpretcast_1357 <= 0;
      __delay_data_2680_plus_1634 <= 0;
      __delay_data_2682_reinterpretcast_1235 <= 0;
      __delay_data_2685__delay_2684_reinterpretcast_1361 <= 0;
      __delay_data_2687_plus_1823 <= 0;
      __delay_data_2689_reinterpretcast_1239 <= 0;
      __delay_data_2692__delay_2691_pointer_1566 <= 0;
      __delay_data_2695__delay_2694_reinterpretcast_1365 <= 0;
      __delay_data_2697_plus_1653 <= 0;
      __delay_data_2699_reinterpretcast_1243 <= 0;
      __delay_data_2702__delay_2701_reinterpretcast_1369 <= 0;
      __delay_data_2704_plus_1842 <= 0;
      __delay_data_2706_reinterpretcast_1247 <= 0;
      __delay_data_2709__delay_2708_pointer_1568 <= 0;
      __delay_data_2712__delay_2711_reinterpretcast_1373 <= 0;
      __delay_data_2714_plus_1672 <= 0;
      __delay_data_2716_reinterpretcast_1251 <= 0;
      __delay_data_2719__delay_2718_reinterpretcast_1377 <= 0;
      __delay_data_2721_plus_1861 <= 0;
      __delay_data_2723_reinterpretcast_1255 <= 0;
      __delay_data_2726__delay_2725_pointer_1570 <= 0;
      __delay_data_2729__delay_2728_reinterpretcast_1381 <= 0;
      __delay_data_2731_plus_1691 <= 0;
      __delay_data_2733_reinterpretcast_1259 <= 0;
      __delay_data_2736__delay_2735_reinterpretcast_1385 <= 0;
      __delay_data_2738_plus_1880 <= 0;
      __delay_data_2740_reinterpretcast_1263 <= 0;
      __delay_data_2743__delay_2742_pointer_1572 <= 0;
      __delay_data_2746__delay_2745_reinterpretcast_1389 <= 0;
      __delay_data_2748_plus_1710 <= 0;
      __delay_data_2750_reinterpretcast_1267 <= 0;
      __delay_data_2753__delay_2752_reinterpretcast_1393 <= 0;
      __delay_data_2755_plus_1899 <= 0;
      __delay_data_2757_reinterpretcast_1271 <= 0;
      __delay_data_2760__delay_2759_pointer_1574 <= 0;
      __delay_data_2763__delay_2762_reinterpretcast_1397 <= 0;
      __delay_data_2765_plus_1729 <= 0;
      __delay_data_2767_reinterpretcast_1275 <= 0;
      __delay_data_2770__delay_2769_reinterpretcast_1401 <= 0;
      __delay_data_2772_plus_1918 <= 0;
      __delay_data_2774_reinterpretcast_1279 <= 0;
      __delay_data_2777__delay_2776_pointer_1576 <= 0;
      __delay_data_2780__delay_2779_reinterpretcast_1405 <= 0;
      __delay_data_2782_plus_1748 <= 0;
      __delay_data_2784_reinterpretcast_1283 <= 0;
      __delay_data_2787__delay_2786_reinterpretcast_1409 <= 0;
      __delay_data_2789_plus_1937 <= 0;
      __delay_data_2791_reinterpretcast_1287 <= 0;
      __delay_data_2794__delay_2793_pointer_1578 <= 0;
      __delay_data_2797__delay_2796_reinterpretcast_1413 <= 0;
      __delay_data_2799_plus_1767 <= 0;
      __delay_data_2801_reinterpretcast_1291 <= 0;
      __delay_data_2804__delay_2803_reinterpretcast_1417 <= 0;
      __delay_data_2806_plus_1956 <= 0;
      __delay_data_2809__delay_2808__variable_951 <= 0;
      __delay_data_2824_plus_1972 <= 0;
      __delay_data_2840__delay_2839__variable_946 <= 0;
      __delay_data_2856__delay_2855_reinterpretcast_1457 <= 0;
      __delay_data_2858_plus_2033 <= 0;
      __delay_data_2861__delay_2860_reinterpretcast_1461 <= 0;
      __delay_data_2863_plus_2222 <= 0;
      __delay_data_2866__delay_2865_reinterpretcast_1465 <= 0;
      __delay_data_2868_plus_2052 <= 0;
      __delay_data_2871__delay_2870_reinterpretcast_1469 <= 0;
      __delay_data_2873_plus_2241 <= 0;
      __delay_data_2876__delay_2875_reinterpretcast_1473 <= 0;
      __delay_data_2878_plus_2071 <= 0;
      __delay_data_2881__delay_2880_reinterpretcast_1477 <= 0;
      __delay_data_2883_plus_2260 <= 0;
      __delay_data_2886__delay_2885_reinterpretcast_1481 <= 0;
      __delay_data_2888_plus_2090 <= 0;
      __delay_data_2891__delay_2890_reinterpretcast_1485 <= 0;
      __delay_data_2893_plus_2279 <= 0;
      __delay_data_2896__delay_2895_reinterpretcast_1489 <= 0;
      __delay_data_2898_plus_2109 <= 0;
      __delay_data_2901__delay_2900_reinterpretcast_1493 <= 0;
      __delay_data_2903_plus_2298 <= 0;
      __delay_data_2906__delay_2905_reinterpretcast_1497 <= 0;
      __delay_data_2908_plus_2128 <= 0;
      __delay_data_2911__delay_2910_reinterpretcast_1501 <= 0;
      __delay_data_2913_plus_2317 <= 0;
      __delay_data_2916__delay_2915_reinterpretcast_1505 <= 0;
      __delay_data_2918_plus_2147 <= 0;
      __delay_data_2921__delay_2920_reinterpretcast_1509 <= 0;
      __delay_data_2923_plus_2336 <= 0;
      __delay_data_2926__delay_2925_reinterpretcast_1513 <= 0;
      __delay_data_2928_plus_2166 <= 0;
      __delay_data_2931__delay_2930_reinterpretcast_1517 <= 0;
      __delay_data_2933_plus_2355 <= 0;
      __delay_data_2936__delay_2935_reinterpretcast_1521 <= 0;
      __delay_data_2938_plus_2185 <= 0;
      __delay_data_2941__delay_2940_reinterpretcast_1525 <= 0;
      __delay_data_2943_plus_2374 <= 0;
      __delay_data_2945_plus_2390 <= 0;
      __delay_data_2961__delay_2960_cond_978 <= 0;
      __delay_data_2983__delay_2982_cond_990 <= 0;
      __delay_data_3005_plus_2409 <= 0;
      __delay_data_3029__delay_3028_cond_977 <= 0;
      __delay_data_3051__delay_3050_cond_989 <= 0;
      __delay_data_3073_plus_1991 <= 0;
      _land_data_960 <= 0;
      _land_data_966 <= 0;
      __delay_data_2654__delay_2653_reinterpretcast_1223 <= 0;
      __delay_data_2657__delay_2656__delay_2655_pointer_1562 <= 0;
      __delay_data_2660__delay_2659__delay_2658_reinterpretcast_1349 <= 0;
      __delay_data_2662__delay_2661_plus_1615 <= 0;
      __delay_data_2666__delay_2665_reinterpretcast_1227 <= 0;
      __delay_data_2669__delay_2668__delay_2667_reinterpretcast_1353 <= 0;
      __delay_data_2671__delay_2670_plus_1804 <= 0;
      __delay_data_2673__delay_2672_reinterpretcast_1231 <= 0;
      __delay_data_2676__delay_2675__delay_2674_pointer_1564 <= 0;
      __delay_data_2679__delay_2678__delay_2677_reinterpretcast_1357 <= 0;
      __delay_data_2681__delay_2680_plus_1634 <= 0;
      __delay_data_2683__delay_2682_reinterpretcast_1235 <= 0;
      __delay_data_2686__delay_2685__delay_2684_reinterpretcast_1361 <= 0;
      __delay_data_2688__delay_2687_plus_1823 <= 0;
      __delay_data_2690__delay_2689_reinterpretcast_1239 <= 0;
      __delay_data_2693__delay_2692__delay_2691_pointer_1566 <= 0;
      __delay_data_2696__delay_2695__delay_2694_reinterpretcast_1365 <= 0;
      __delay_data_2698__delay_2697_plus_1653 <= 0;
      __delay_data_2700__delay_2699_reinterpretcast_1243 <= 0;
      __delay_data_2703__delay_2702__delay_2701_reinterpretcast_1369 <= 0;
      __delay_data_2705__delay_2704_plus_1842 <= 0;
      __delay_data_2707__delay_2706_reinterpretcast_1247 <= 0;
      __delay_data_2710__delay_2709__delay_2708_pointer_1568 <= 0;
      __delay_data_2713__delay_2712__delay_2711_reinterpretcast_1373 <= 0;
      __delay_data_2715__delay_2714_plus_1672 <= 0;
      __delay_data_2717__delay_2716_reinterpretcast_1251 <= 0;
      __delay_data_2720__delay_2719__delay_2718_reinterpretcast_1377 <= 0;
      __delay_data_2722__delay_2721_plus_1861 <= 0;
      __delay_data_2724__delay_2723_reinterpretcast_1255 <= 0;
      __delay_data_2727__delay_2726__delay_2725_pointer_1570 <= 0;
      __delay_data_2730__delay_2729__delay_2728_reinterpretcast_1381 <= 0;
      __delay_data_2732__delay_2731_plus_1691 <= 0;
      __delay_data_2734__delay_2733_reinterpretcast_1259 <= 0;
      __delay_data_2737__delay_2736__delay_2735_reinterpretcast_1385 <= 0;
      __delay_data_2739__delay_2738_plus_1880 <= 0;
      __delay_data_2741__delay_2740_reinterpretcast_1263 <= 0;
      __delay_data_2744__delay_2743__delay_2742_pointer_1572 <= 0;
      __delay_data_2747__delay_2746__delay_2745_reinterpretcast_1389 <= 0;
      __delay_data_2749__delay_2748_plus_1710 <= 0;
      __delay_data_2751__delay_2750_reinterpretcast_1267 <= 0;
      __delay_data_2754__delay_2753__delay_2752_reinterpretcast_1393 <= 0;
      __delay_data_2756__delay_2755_plus_1899 <= 0;
      __delay_data_2758__delay_2757_reinterpretcast_1271 <= 0;
      __delay_data_2761__delay_2760__delay_2759_pointer_1574 <= 0;
      __delay_data_2764__delay_2763__delay_2762_reinterpretcast_1397 <= 0;
      __delay_data_2766__delay_2765_plus_1729 <= 0;
      __delay_data_2768__delay_2767_reinterpretcast_1275 <= 0;
      __delay_data_2771__delay_2770__delay_2769_reinterpretcast_1401 <= 0;
      __delay_data_2773__delay_2772_plus_1918 <= 0;
      __delay_data_2775__delay_2774_reinterpretcast_1279 <= 0;
      __delay_data_2778__delay_2777__delay_2776_pointer_1576 <= 0;
      __delay_data_2781__delay_2780__delay_2779_reinterpretcast_1405 <= 0;
      __delay_data_2783__delay_2782_plus_1748 <= 0;
      __delay_data_2785__delay_2784_reinterpretcast_1283 <= 0;
      __delay_data_2788__delay_2787__delay_2786_reinterpretcast_1409 <= 0;
      __delay_data_2790__delay_2789_plus_1937 <= 0;
      __delay_data_2792__delay_2791_reinterpretcast_1287 <= 0;
      __delay_data_2795__delay_2794__delay_2793_pointer_1578 <= 0;
      __delay_data_2798__delay_2797__delay_2796_reinterpretcast_1413 <= 0;
      __delay_data_2800__delay_2799_plus_1767 <= 0;
      __delay_data_2802__delay_2801_reinterpretcast_1291 <= 0;
      __delay_data_2805__delay_2804__delay_2803_reinterpretcast_1417 <= 0;
      __delay_data_2807__delay_2806_plus_1956 <= 0;
      __delay_data_2810__delay_2809__delay_2808__variable_951 <= 0;
      __delay_data_2825__delay_2824_plus_1972 <= 0;
      __delay_data_2841__delay_2840__delay_2839__variable_946 <= 0;
      __delay_data_2857__delay_2856__delay_2855_reinterpretcast_1457 <= 0;
      __delay_data_2859__delay_2858_plus_2033 <= 0;
      __delay_data_2862__delay_2861__delay_2860_reinterpretcast_1461 <= 0;
      __delay_data_2864__delay_2863_plus_2222 <= 0;
      __delay_data_2867__delay_2866__delay_2865_reinterpretcast_1465 <= 0;
      __delay_data_2869__delay_2868_plus_2052 <= 0;
      __delay_data_2872__delay_2871__delay_2870_reinterpretcast_1469 <= 0;
      __delay_data_2874__delay_2873_plus_2241 <= 0;
      __delay_data_2877__delay_2876__delay_2875_reinterpretcast_1473 <= 0;
      __delay_data_2879__delay_2878_plus_2071 <= 0;
      __delay_data_2882__delay_2881__delay_2880_reinterpretcast_1477 <= 0;
      __delay_data_2884__delay_2883_plus_2260 <= 0;
      __delay_data_2887__delay_2886__delay_2885_reinterpretcast_1481 <= 0;
      __delay_data_2889__delay_2888_plus_2090 <= 0;
      __delay_data_2892__delay_2891__delay_2890_reinterpretcast_1485 <= 0;
      __delay_data_2894__delay_2893_plus_2279 <= 0;
      __delay_data_2897__delay_2896__delay_2895_reinterpretcast_1489 <= 0;
      __delay_data_2899__delay_2898_plus_2109 <= 0;
      __delay_data_2902__delay_2901__delay_2900_reinterpretcast_1493 <= 0;
      __delay_data_2904__delay_2903_plus_2298 <= 0;
      __delay_data_2907__delay_2906__delay_2905_reinterpretcast_1497 <= 0;
      __delay_data_2909__delay_2908_plus_2128 <= 0;
      __delay_data_2912__delay_2911__delay_2910_reinterpretcast_1501 <= 0;
      __delay_data_2914__delay_2913_plus_2317 <= 0;
      __delay_data_2917__delay_2916__delay_2915_reinterpretcast_1505 <= 0;
      __delay_data_2919__delay_2918_plus_2147 <= 0;
      __delay_data_2922__delay_2921__delay_2920_reinterpretcast_1509 <= 0;
      __delay_data_2924__delay_2923_plus_2336 <= 0;
      __delay_data_2927__delay_2926__delay_2925_reinterpretcast_1513 <= 0;
      __delay_data_2929__delay_2928_plus_2166 <= 0;
      __delay_data_2932__delay_2931__delay_2930_reinterpretcast_1517 <= 0;
      __delay_data_2934__delay_2933_plus_2355 <= 0;
      __delay_data_2937__delay_2936__delay_2935_reinterpretcast_1521 <= 0;
      __delay_data_2939__delay_2938_plus_2185 <= 0;
      __delay_data_2942__delay_2941__delay_2940_reinterpretcast_1525 <= 0;
      __delay_data_2944__delay_2943_plus_2374 <= 0;
      __delay_data_2946__delay_2945_plus_2390 <= 0;
      __delay_data_2962__delay_2961__delay_2960_cond_978 <= 0;
      __delay_data_2984__delay_2983__delay_2982_cond_990 <= 0;
      __delay_data_3006__delay_3005_plus_2409 <= 0;
      __delay_data_3030__delay_3029__delay_3028_cond_977 <= 0;
      __delay_data_3052__delay_3051__delay_3050_cond_989 <= 0;
      __delay_data_3074__delay_3073_plus_1991 <= 0;
      __delay_data_2811__delay_2810__delay_2809____variable_951 <= 0;
      __delay_data_2826__delay_2825__delay_2824_plus_1972 <= 0;
      __delay_data_2842__delay_2841__delay_2840____variable_946 <= 0;
      __delay_data_2947__delay_2946__delay_2945_plus_2390 <= 0;
      __delay_data_2963__delay_2962__delay_2961__delay_2960_cond_978 <= 0;
      __delay_data_2985__delay_2984__delay_2983__delay_2982_cond_990 <= 0;
      __delay_data_3007__delay_3006__delay_3005_plus_2409 <= 0;
      __delay_data_3031__delay_3030__delay_3029__delay_3028_cond_977 <= 0;
      __delay_data_3053__delay_3052__delay_3051__delay_3050_cond_989 <= 0;
      __delay_data_3075__delay_3074__delay_3073_plus_1991 <= 0;
      __delay_data_2812__delay_2811__delay_2810____variable_951 <= 0;
      __delay_data_2827__delay_2826__delay_2825___plus_1972 <= 0;
      __delay_data_2843__delay_2842__delay_2841____variable_946 <= 0;
      __delay_data_2948__delay_2947__delay_2946___plus_2390 <= 0;
      __delay_data_2964__delay_2963__delay_2962__delay_2961___cond_978 <= 0;
      __delay_data_2986__delay_2985__delay_2984__delay_2983___cond_990 <= 0;
      __delay_data_3008__delay_3007__delay_3006___plus_2409 <= 0;
      __delay_data_3032__delay_3031__delay_3030__delay_3029___cond_977 <= 0;
      __delay_data_3054__delay_3053__delay_3052__delay_3051___cond_989 <= 0;
      __delay_data_3076__delay_3075__delay_3074___plus_1991 <= 0;
      __delay_data_2813__delay_2812__delay_2811____variable_951 <= 0;
      __delay_data_2828__delay_2827__delay_2826___plus_1972 <= 0;
      __delay_data_2844__delay_2843__delay_2842____variable_946 <= 0;
      __delay_data_2949__delay_2948__delay_2947___plus_2390 <= 0;
      __delay_data_2965__delay_2964__delay_2963__delay_2962___cond_978 <= 0;
      __delay_data_2987__delay_2986__delay_2985__delay_2984___cond_990 <= 0;
      __delay_data_3009__delay_3008__delay_3007___plus_2409 <= 0;
      __delay_data_3033__delay_3032__delay_3031__delay_3030___cond_977 <= 0;
      __delay_data_3055__delay_3054__delay_3053__delay_3052___cond_989 <= 0;
      __delay_data_3077__delay_3076__delay_3075___plus_1991 <= 0;
      __delay_data_2814__delay_2813__delay_2812____variable_951 <= 0;
      __delay_data_2829__delay_2828__delay_2827___plus_1972 <= 0;
      __delay_data_2845__delay_2844__delay_2843____variable_946 <= 0;
      __delay_data_2950__delay_2949__delay_2948___plus_2390 <= 0;
      __delay_data_2966__delay_2965__delay_2964__delay_2963___cond_978 <= 0;
      __delay_data_2988__delay_2987__delay_2986__delay_2985___cond_990 <= 0;
      __delay_data_3010__delay_3009__delay_3008___plus_2409 <= 0;
      __delay_data_3034__delay_3033__delay_3032__delay_3031___cond_977 <= 0;
      __delay_data_3056__delay_3055__delay_3054__delay_3053___cond_989 <= 0;
      __delay_data_3078__delay_3077__delay_3076___plus_1991 <= 0;
      __delay_data_2815__delay_2814__delay_2813____variable_951 <= 0;
      __delay_data_2830__delay_2829__delay_2828___plus_1972 <= 0;
      __delay_data_2846__delay_2845__delay_2844____variable_946 <= 0;
      __delay_data_2951__delay_2950__delay_2949___plus_2390 <= 0;
      __delay_data_2967__delay_2966__delay_2965__delay_2964___cond_978 <= 0;
      __delay_data_2989__delay_2988__delay_2987__delay_2986___cond_990 <= 0;
      __delay_data_3011__delay_3010__delay_3009___plus_2409 <= 0;
      __delay_data_3035__delay_3034__delay_3033__delay_3032___cond_977 <= 0;
      __delay_data_3057__delay_3056__delay_3055__delay_3054___cond_989 <= 0;
      __delay_data_3079__delay_3078__delay_3077___plus_1991 <= 0;
      __delay_data_2816__delay_2815__delay_2814____variable_951 <= 0;
      __delay_data_2831__delay_2830__delay_2829___plus_1972 <= 0;
      __delay_data_2847__delay_2846__delay_2845____variable_946 <= 0;
      __delay_data_2952__delay_2951__delay_2950___plus_2390 <= 0;
      __delay_data_2968__delay_2967__delay_2966__delay_2965___cond_978 <= 0;
      __delay_data_2990__delay_2989__delay_2988__delay_2987___cond_990 <= 0;
      __delay_data_3012__delay_3011__delay_3010___plus_2409 <= 0;
      __delay_data_3036__delay_3035__delay_3034__delay_3033___cond_977 <= 0;
      __delay_data_3058__delay_3057__delay_3056__delay_3055___cond_989 <= 0;
      __delay_data_3080__delay_3079__delay_3078___plus_1991 <= 0;
      __delay_data_2817__delay_2816__delay_2815____variable_951 <= 0;
      __delay_data_2832__delay_2831__delay_2830___plus_1972 <= 0;
      __delay_data_2848__delay_2847__delay_2846____variable_946 <= 0;
      __delay_data_2953__delay_2952__delay_2951___plus_2390 <= 0;
      __delay_data_2969__delay_2968__delay_2967__delay_2966___cond_978 <= 0;
      __delay_data_2991__delay_2990__delay_2989__delay_2988___cond_990 <= 0;
      __delay_data_3013__delay_3012__delay_3011___plus_2409 <= 0;
      __delay_data_3037__delay_3036__delay_3035__delay_3034___cond_977 <= 0;
      __delay_data_3059__delay_3058__delay_3057__delay_3056___cond_989 <= 0;
      __delay_data_3081__delay_3080__delay_3079___plus_1991 <= 0;
      __delay_data_2818__delay_2817__delay_2816____variable_951 <= 0;
      __delay_data_2833__delay_2832__delay_2831___plus_1972 <= 0;
      __delay_data_2849__delay_2848__delay_2847____variable_946 <= 0;
      __delay_data_2954__delay_2953__delay_2952___plus_2390 <= 0;
      __delay_data_2970__delay_2969__delay_2968__delay_2967___cond_978 <= 0;
      __delay_data_2992__delay_2991__delay_2990__delay_2989___cond_990 <= 0;
      __delay_data_3014__delay_3013__delay_3012___plus_2409 <= 0;
      __delay_data_3038__delay_3037__delay_3036__delay_3035___cond_977 <= 0;
      __delay_data_3060__delay_3059__delay_3058__delay_3057___cond_989 <= 0;
      __delay_data_3082__delay_3081__delay_3080___plus_1991 <= 0;
      __delay_data_2819__delay_2818__delay_2817____variable_951 <= 0;
      __delay_data_2834__delay_2833__delay_2832___plus_1972 <= 0;
      __delay_data_2850__delay_2849__delay_2848____variable_946 <= 0;
      __delay_data_2955__delay_2954__delay_2953___plus_2390 <= 0;
      __delay_data_2971__delay_2970__delay_2969__delay_2968___cond_978 <= 0;
      __delay_data_2993__delay_2992__delay_2991__delay_2990___cond_990 <= 0;
      __delay_data_3015__delay_3014__delay_3013___plus_2409 <= 0;
      __delay_data_3039__delay_3038__delay_3037__delay_3036___cond_977 <= 0;
      __delay_data_3061__delay_3060__delay_3059__delay_3058___cond_989 <= 0;
      __delay_data_3083__delay_3082__delay_3081___plus_1991 <= 0;
      __delay_data_2820__delay_2819__delay_2818____variable_951 <= 0;
      __delay_data_2835__delay_2834__delay_2833___plus_1972 <= 0;
      __delay_data_2851__delay_2850__delay_2849____variable_946 <= 0;
      __delay_data_2956__delay_2955__delay_2954___plus_2390 <= 0;
      __delay_data_2972__delay_2971__delay_2970__delay_2969___cond_978 <= 0;
      __delay_data_2994__delay_2993__delay_2992__delay_2991___cond_990 <= 0;
      __delay_data_3016__delay_3015__delay_3014___plus_2409 <= 0;
      __delay_data_3040__delay_3039__delay_3038__delay_3037___cond_977 <= 0;
      __delay_data_3062__delay_3061__delay_3060__delay_3059___cond_989 <= 0;
      __delay_data_3084__delay_3083__delay_3082___plus_1991 <= 0;
      __delay_data_2821__delay_2820__delay_2819____variable_951 <= 0;
      __delay_data_2836__delay_2835__delay_2834___plus_1972 <= 0;
      __delay_data_2852__delay_2851__delay_2850____variable_946 <= 0;
      __delay_data_2957__delay_2956__delay_2955___plus_2390 <= 0;
      __delay_data_2973__delay_2972__delay_2971__delay_2970___cond_978 <= 0;
      __delay_data_2995__delay_2994__delay_2993__delay_2992___cond_990 <= 0;
      __delay_data_3017__delay_3016__delay_3015___plus_2409 <= 0;
      __delay_data_3041__delay_3040__delay_3039__delay_3038___cond_977 <= 0;
      __delay_data_3063__delay_3062__delay_3061__delay_3060___cond_989 <= 0;
      __delay_data_3085__delay_3084__delay_3083___plus_1991 <= 0;
      __delay_data_2822__delay_2821__delay_2820____variable_951 <= 0;
      __delay_data_2837__delay_2836__delay_2835___plus_1972 <= 0;
      __delay_data_2853__delay_2852__delay_2851____variable_946 <= 0;
      __delay_data_2958__delay_2957__delay_2956___plus_2390 <= 0;
      __delay_data_2974__delay_2973__delay_2972__delay_2971___cond_978 <= 0;
      __delay_data_2996__delay_2995__delay_2994__delay_2993___cond_990 <= 0;
      __delay_data_3018__delay_3017__delay_3016___plus_2409 <= 0;
      __delay_data_3042__delay_3041__delay_3040__delay_3039___cond_977 <= 0;
      __delay_data_3064__delay_3063__delay_3062__delay_3061___cond_989 <= 0;
      __delay_data_3086__delay_3085__delay_3084___plus_1991 <= 0;
      __delay_data_2823__delay_2822__delay_2821____variable_951 <= 0;
      __delay_data_2838__delay_2837__delay_2836___plus_1972 <= 0;
      __delay_data_2854__delay_2853__delay_2852____variable_946 <= 0;
      __delay_data_2959__delay_2958__delay_2957___plus_2390 <= 0;
      __delay_data_2975__delay_2974__delay_2973__delay_2972___cond_978 <= 0;
      __delay_data_2997__delay_2996__delay_2995__delay_2994___cond_990 <= 0;
      __delay_data_3019__delay_3018__delay_3017___plus_2409 <= 0;
      __delay_data_3043__delay_3042__delay_3041__delay_3040___cond_977 <= 0;
      __delay_data_3065__delay_3064__delay_3063__delay_3062___cond_989 <= 0;
      __delay_data_3087__delay_3086__delay_3085___plus_1991 <= 0;
      __delay_data_2976__delay_2975__delay_2974__delay_2973___cond_978 <= 0;
      __delay_data_2998__delay_2997__delay_2996__delay_2995___cond_990 <= 0;
      __delay_data_3020__delay_3019__delay_3018___plus_2409 <= 0;
      __delay_data_3044__delay_3043__delay_3042__delay_3041___cond_977 <= 0;
      __delay_data_3066__delay_3065__delay_3064__delay_3063___cond_989 <= 0;
      __delay_data_3088__delay_3087__delay_3086___plus_1991 <= 0;
      __delay_data_2977__delay_2976__delay_2975__delay_2974___cond_978 <= 0;
      __delay_data_2999__delay_2998__delay_2997__delay_2996___cond_990 <= 0;
      __delay_data_3021__delay_3020__delay_3019___plus_2409 <= 0;
      __delay_data_3045__delay_3044__delay_3043__delay_3042___cond_977 <= 0;
      __delay_data_3067__delay_3066__delay_3065__delay_3064___cond_989 <= 0;
      __delay_data_3089__delay_3088__delay_3087___plus_1991 <= 0;
      __delay_data_2978__delay_2977__delay_2976__delay_2975___cond_978 <= 0;
      __delay_data_3000__delay_2999__delay_2998__delay_2997___cond_990 <= 0;
      __delay_data_3022__delay_3021__delay_3020___plus_2409 <= 0;
      __delay_data_3046__delay_3045__delay_3044__delay_3043___cond_977 <= 0;
      __delay_data_3068__delay_3067__delay_3066__delay_3065___cond_989 <= 0;
      __delay_data_3090__delay_3089__delay_3088___plus_1991 <= 0;
      __delay_data_2979__delay_2978__delay_2977__delay_2976___cond_978 <= 0;
      __delay_data_3001__delay_3000__delay_2999__delay_2998___cond_990 <= 0;
      __delay_data_3023__delay_3022__delay_3021___plus_2409 <= 0;
      __delay_data_3047__delay_3046__delay_3045__delay_3044___cond_977 <= 0;
      __delay_data_3069__delay_3068__delay_3067__delay_3066___cond_989 <= 0;
      __delay_data_3091__delay_3090__delay_3089___plus_1991 <= 0;
      __delay_data_2980__delay_2979__delay_2978__delay_2977___cond_978 <= 0;
      __delay_data_3002__delay_3001__delay_3000__delay_2999___cond_990 <= 0;
      __delay_data_3024__delay_3023__delay_3022___plus_2409 <= 0;
      __delay_data_3048__delay_3047__delay_3046__delay_3045___cond_977 <= 0;
      __delay_data_3070__delay_3069__delay_3068__delay_3067___cond_989 <= 0;
      __delay_data_3092__delay_3091__delay_3090___plus_1991 <= 0;
      __delay_data_2981__delay_2980__delay_2979__delay_2978___cond_978 <= 0;
      __delay_data_3003__delay_3002__delay_3001__delay_3000___cond_990 <= 0;
      __delay_data_3025__delay_3024__delay_3023___plus_2409 <= 0;
      __delay_data_3049__delay_3048__delay_3047__delay_3046___cond_977 <= 0;
      __delay_data_3071__delay_3070__delay_3069__delay_3068___cond_989 <= 0;
      __delay_data_3093__delay_3092__delay_3091___plus_1991 <= 0;
      _plus_data_1975 <= 0;
      _plus_data_2393 <= 0;
      __delay_data_3004__delay_3003__delay_3002__delay_3001___cond_990 <= 0;
      __delay_data_3026__delay_3025__delay_3024___plus_2409 <= 0;
      __delay_data_3072__delay_3071__delay_3070__delay_3069___cond_989 <= 0;
      __delay_data_3094__delay_3093__delay_3092___plus_1991 <= 0;
      __delay_data_3096__substreamoutput_1974 <= 0;
      __delay_data_3097__delay_3096__substreamoutput_1974 <= 0;
      __delay_data_3098__delay_3097____substreamoutput_1974 <= 0;
      __delay_data_3099__delay_3098____substreamoutput_1974 <= 0;
      __delay_data_3100__delay_3099____substreamoutput_1974 <= 0;
      __delay_data_3101__delay_3100____substreamoutput_1974 <= 0;
      __delay_data_3102__delay_3101____substreamoutput_1974 <= 0;
      __delay_data_3103__delay_3102____substreamoutput_1974 <= 0;
      __delay_data_3104__delay_3103____substreamoutput_1974 <= 0;
      __delay_data_3105__delay_3104____substreamoutput_1974 <= 0;
      _greaterthan_data_1994 <= 0;
      _greaterthan_data_2412 <= 0;
      __delay_data_3027__substreamoutput_2410 <= 0;
      __delay_data_3095__substreamoutput_1992 <= 0;
      __delay_data_3106__delay_3105____substreamoutput_1974 <= 0;
      _cond_data_1996 <= 0;
      _cond_data_2414 <= 0;
      __delay_data_3107__delay_3106____substreamoutput_1974 <= 0;
      _stream_conv2d_4_parameter_0_next_parameter_data <= 0;
      __variable_wdata_946 <= 0;
      _stream_conv2d_4_parameter_1_next_parameter_data <= 0;
      __variable_wdata_947 <= 0;
      _stream_conv2d_4_parameter_2_next_parameter_data <= 0;
      __variable_wdata_948 <= 0;
      _stream_conv2d_4_parameter_3_next_parameter_data <= 0;
      __variable_wdata_949 <= 0;
      _stream_conv2d_4_parameter_4_next_parameter_data <= 0;
      __variable_wdata_950 <= 0;
      _stream_conv2d_4_parameter_6_next_parameter_data <= 0;
      __variable_wdata_967 <= 0;
      _stream_conv2d_4_source_7_source_mode <= 5'b0;
      _stream_conv2d_4_source_7_source_offset <= 0;
      _source_stream_conv2d_4_source_7_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_3 <= 0;
      _stream_conv2d_4_source_7_source_sel <= 0;
      _stream_conv2d_4_source_7_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_968 <= 0;
      _stream_conv2d_4_source_7_source_ram_raddr <= 0;
      _stream_conv2d_4_parameter_8_next_parameter_data <= 0;
      __variable_wdata_979 <= 0;
      _stream_conv2d_4_source_9_source_mode <= 5'b0;
      _stream_conv2d_4_source_9_source_offset <= 0;
      _source_stream_conv2d_4_source_9_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_3 <= 0;
      _stream_conv2d_4_source_9_source_sel <= 0;
      _stream_conv2d_4_source_9_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_980 <= 0;
      _stream_conv2d_4_source_9_source_ram_raddr <= 0;
      _stream_conv2d_4_parameter_10_next_parameter_data <= 0;
      __variable_wdata_991 <= 0;
      _stream_conv2d_4_source_11_source_mode <= 5'b0;
      _stream_conv2d_4_source_11_source_empty_data <= 0;
      __variable_wdata_992 <= 0;
      _stream_conv2d_4_parameter_12_next_parameter_data <= 0;
      __variable_wdata_1003 <= 0;
      _stream_conv2d_4_source_13_source_mode <= 5'b0;
      _stream_conv2d_4_source_13_source_empty_data <= 0;
      __variable_wdata_1004 <= 0;
      _stream_conv2d_4_parameter_14_next_parameter_data <= 0;
      __variable_wdata_1015 <= 0;
      _stream_conv2d_4_source_15_source_mode <= 5'b0;
      _stream_conv2d_4_source_15_source_empty_data <= 0;
      __variable_wdata_1016 <= 0;
      _stream_conv2d_4_parameter_16_next_parameter_data <= 0;
      __variable_wdata_1027 <= 0;
      _stream_conv2d_4_parameter_17_next_parameter_data <= 0;
      __variable_wdata_1028 <= 0;
      _stream_conv2d_4_parameter_18_next_parameter_data <= 0;
      __variable_wdata_1029 <= 0;
      _stream_conv2d_4_parameter_19_next_parameter_data <= 0;
      __variable_wdata_1030 <= 0;
      _stream_conv2d_4_source_20_source_mode <= 5'b0;
      _stream_conv2d_4_source_20_source_offset <= 0;
      _source_stream_conv2d_4_source_20_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_3 <= 0;
      _stream_conv2d_4_source_20_source_sel <= 0;
      _stream_conv2d_4_source_20_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_1031 <= 0;
      _stream_conv2d_4_source_20_source_ram_raddr <= 0;
      _stream_conv2d_4_source_21_source_mode <= 5'b0;
      _stream_conv2d_4_source_21_source_offset <= 0;
      _source_stream_conv2d_4_source_21_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_3 <= 0;
      _stream_conv2d_4_source_21_source_sel <= 0;
      _stream_conv2d_4_source_21_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_1032 <= 0;
      _stream_conv2d_4_source_21_source_ram_raddr <= 0;
      _stream_conv2d_4_source_22_source_mode <= 5'b0;
      _stream_conv2d_4_source_22_source_offset <= 0;
      _source_stream_conv2d_4_source_22_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_3 <= 0;
      _stream_conv2d_4_source_22_source_sel <= 0;
      _stream_conv2d_4_source_22_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_1033 <= 0;
      _stream_conv2d_4_source_22_source_ram_raddr <= 0;
      _stream_conv2d_4_source_23_source_mode <= 5'b0;
      _stream_conv2d_4_source_23_source_offset <= 0;
      _source_stream_conv2d_4_source_23_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_3 <= 0;
      _stream_conv2d_4_source_23_source_sel <= 0;
      _stream_conv2d_4_source_23_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_3 <= 0;
      __variable_wdata_1034 <= 0;
      _stream_conv2d_4_source_23_source_ram_raddr <= 0;
      _stream_conv2d_4_source_24_source_mode <= 5'b0;
      _stream_conv2d_4_source_24_source_offset <= 0;
      _source_stream_conv2d_4_source_24_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_3 <= 0;
      _stream_conv2d_4_source_24_source_sel <= 0;
      _stream_conv2d_4_source_24_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_3 <= 0;
      __variable_wdata_1035 <= 0;
      _stream_conv2d_4_source_24_source_ram_raddr <= 0;
      _stream_conv2d_4_source_25_source_mode <= 5'b0;
      _stream_conv2d_4_source_25_source_offset <= 0;
      _source_stream_conv2d_4_source_25_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_3 <= 0;
      _stream_conv2d_4_source_25_source_sel <= 0;
      _stream_conv2d_4_source_25_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_3 <= 0;
      __variable_wdata_1036 <= 0;
      _stream_conv2d_4_source_25_source_ram_raddr <= 0;
      _stream_conv2d_4_source_26_source_mode <= 5'b0;
      _stream_conv2d_4_source_26_source_offset <= 0;
      _source_stream_conv2d_4_source_26_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_3 <= 0;
      _stream_conv2d_4_source_26_source_sel <= 0;
      _stream_conv2d_4_source_26_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_3 <= 0;
      __variable_wdata_1037 <= 0;
      _stream_conv2d_4_source_26_source_ram_raddr <= 0;
      _stream_conv2d_4_source_27_source_mode <= 5'b0;
      _stream_conv2d_4_source_27_source_offset <= 0;
      _source_stream_conv2d_4_source_27_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_3 <= 0;
      _stream_conv2d_4_source_27_source_sel <= 0;
      _stream_conv2d_4_source_27_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_3 <= 0;
      __variable_wdata_1038 <= 0;
      _stream_conv2d_4_source_27_source_ram_raddr <= 0;
      _stream_conv2d_4_source_28_source_mode <= 5'b0;
      _stream_conv2d_4_source_28_source_offset <= 0;
      _source_stream_conv2d_4_source_28_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_3 <= 0;
      _stream_conv2d_4_source_28_source_sel <= 0;
      _stream_conv2d_4_source_28_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_3 <= 0;
      __variable_wdata_1039 <= 0;
      _stream_conv2d_4_source_28_source_ram_raddr <= 0;
      _stream_conv2d_4_source_29_source_mode <= 5'b0;
      _stream_conv2d_4_source_29_source_offset <= 0;
      _source_stream_conv2d_4_source_29_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_3 <= 0;
      _stream_conv2d_4_source_29_source_sel <= 0;
      _stream_conv2d_4_source_29_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_3 <= 0;
      __variable_wdata_1328 <= 0;
      _stream_conv2d_4_source_29_source_ram_raddr <= 0;
      _stream_conv2d_4_source_30_source_mode <= 5'b0;
      _stream_conv2d_4_source_30_source_offset <= 0;
      _source_stream_conv2d_4_source_30_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_3 <= 0;
      _stream_conv2d_4_source_30_source_sel <= 0;
      _stream_conv2d_4_source_30_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_3 <= 0;
      __variable_wdata_1329 <= 0;
      _stream_conv2d_4_source_30_source_ram_raddr <= 0;
      _stream_conv2d_4_source_31_source_mode <= 5'b0;
      _stream_conv2d_4_source_31_source_offset <= 0;
      _source_stream_conv2d_4_source_31_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_3 <= 0;
      _stream_conv2d_4_source_31_source_sel <= 0;
      _stream_conv2d_4_source_31_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_3 <= 0;
      __variable_wdata_1330 <= 0;
      _stream_conv2d_4_source_31_source_ram_raddr <= 0;
      _stream_conv2d_4_source_32_source_mode <= 5'b0;
      _stream_conv2d_4_source_32_source_offset <= 0;
      _source_stream_conv2d_4_source_32_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_3 <= 0;
      _stream_conv2d_4_source_32_source_sel <= 0;
      _stream_conv2d_4_source_32_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_3 <= 0;
      __variable_wdata_1331 <= 0;
      _stream_conv2d_4_source_32_source_ram_raddr <= 0;
      _stream_conv2d_4_source_33_source_mode <= 5'b0;
      _stream_conv2d_4_source_33_source_offset <= 0;
      _source_stream_conv2d_4_source_33_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_3 <= 0;
      _stream_conv2d_4_source_33_source_sel <= 0;
      _stream_conv2d_4_source_33_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_3 <= 0;
      __variable_wdata_1332 <= 0;
      _stream_conv2d_4_source_33_source_ram_raddr <= 0;
      _stream_conv2d_4_source_34_source_mode <= 5'b0;
      _stream_conv2d_4_source_34_source_offset <= 0;
      _source_stream_conv2d_4_source_34_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_3 <= 0;
      _stream_conv2d_4_source_34_source_sel <= 0;
      _stream_conv2d_4_source_34_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_3 <= 0;
      __variable_wdata_1333 <= 0;
      _stream_conv2d_4_source_34_source_ram_raddr <= 0;
      _stream_conv2d_4_source_35_source_mode <= 5'b0;
      _stream_conv2d_4_source_35_source_offset <= 0;
      _source_stream_conv2d_4_source_35_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_3 <= 0;
      _stream_conv2d_4_source_35_source_sel <= 0;
      _stream_conv2d_4_source_35_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_3 <= 0;
      __variable_wdata_1334 <= 0;
      _stream_conv2d_4_source_35_source_ram_raddr <= 0;
      _stream_conv2d_4_source_36_source_mode <= 5'b0;
      _stream_conv2d_4_source_36_source_offset <= 0;
      _source_stream_conv2d_4_source_36_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_3 <= 0;
      _stream_conv2d_4_source_36_source_sel <= 0;
      _stream_conv2d_4_source_36_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_3 <= 0;
      __variable_wdata_1335 <= 0;
      _stream_conv2d_4_source_36_source_ram_raddr <= 0;
      _stream_conv2d_4_source_37_source_mode <= 5'b0;
      _stream_conv2d_4_source_37_source_offset <= 0;
      _source_stream_conv2d_4_source_37_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_3 <= 0;
      _stream_conv2d_4_source_37_source_sel <= 0;
      _stream_conv2d_4_source_37_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_3 <= 0;
      __variable_wdata_1336 <= 0;
      _stream_conv2d_4_source_37_source_ram_raddr <= 0;
      _stream_conv2d_4_source_38_source_mode <= 5'b0;
      _stream_conv2d_4_source_38_source_offset <= 0;
      _source_stream_conv2d_4_source_38_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_38_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_38_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_38_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_3 <= 0;
      _stream_conv2d_4_source_38_source_sel <= 0;
      _stream_conv2d_4_source_38_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_38_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_38_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_38_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_38_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_38_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_38_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_38_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_38_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_38_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_38_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_38_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_38_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_38_pat_stride_buf_3 <= 0;
      __variable_wdata_1337 <= 0;
      _stream_conv2d_4_source_38_source_ram_raddr <= 0;
      _stream_conv2d_4_source_39_source_mode <= 5'b0;
      _stream_conv2d_4_source_39_source_offset <= 0;
      _source_stream_conv2d_4_source_39_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_39_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_39_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_39_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_3 <= 0;
      _stream_conv2d_4_source_39_source_sel <= 0;
      _stream_conv2d_4_source_39_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_39_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_39_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_39_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_39_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_39_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_39_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_39_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_39_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_39_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_39_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_39_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_39_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_39_pat_stride_buf_3 <= 0;
      __variable_wdata_1338 <= 0;
      _stream_conv2d_4_source_39_source_ram_raddr <= 0;
      _stream_conv2d_4_source_40_source_mode <= 5'b0;
      _stream_conv2d_4_source_40_source_offset <= 0;
      _source_stream_conv2d_4_source_40_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_40_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_40_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_40_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_3 <= 0;
      _stream_conv2d_4_source_40_source_sel <= 0;
      _stream_conv2d_4_source_40_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_40_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_40_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_40_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_40_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_40_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_40_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_40_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_40_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_40_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_40_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_40_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_40_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_40_pat_stride_buf_3 <= 0;
      __variable_wdata_1339 <= 0;
      _stream_conv2d_4_source_40_source_ram_raddr <= 0;
      _stream_conv2d_4_source_41_source_mode <= 5'b0;
      _stream_conv2d_4_source_41_source_offset <= 0;
      _source_stream_conv2d_4_source_41_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_41_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_41_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_41_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_3 <= 0;
      _stream_conv2d_4_source_41_source_sel <= 0;
      _stream_conv2d_4_source_41_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_41_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_41_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_41_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_41_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_41_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_41_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_41_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_41_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_41_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_41_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_41_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_41_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_41_pat_stride_buf_3 <= 0;
      __variable_wdata_1340 <= 0;
      _stream_conv2d_4_source_41_source_ram_raddr <= 0;
      _stream_conv2d_4_source_42_source_mode <= 5'b0;
      _stream_conv2d_4_source_42_source_offset <= 0;
      _source_stream_conv2d_4_source_42_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_42_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_42_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_42_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_3 <= 0;
      _stream_conv2d_4_source_42_source_sel <= 0;
      _stream_conv2d_4_source_42_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_42_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_42_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_42_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_42_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_42_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_42_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_42_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_42_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_42_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_42_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_42_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_42_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_42_pat_stride_buf_3 <= 0;
      __variable_wdata_1341 <= 0;
      _stream_conv2d_4_source_42_source_ram_raddr <= 0;
      _stream_conv2d_4_source_43_source_mode <= 5'b0;
      _stream_conv2d_4_source_43_source_offset <= 0;
      _source_stream_conv2d_4_source_43_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_43_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_43_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_43_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_3 <= 0;
      _stream_conv2d_4_source_43_source_sel <= 0;
      _stream_conv2d_4_source_43_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_43_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_43_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_43_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_43_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_43_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_43_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_43_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_43_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_43_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_43_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_43_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_43_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_43_pat_stride_buf_3 <= 0;
      __variable_wdata_1342 <= 0;
      _stream_conv2d_4_source_43_source_ram_raddr <= 0;
      _stream_conv2d_4_source_44_source_mode <= 5'b0;
      _stream_conv2d_4_source_44_source_offset <= 0;
      _source_stream_conv2d_4_source_44_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_44_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_44_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_44_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_3 <= 0;
      _stream_conv2d_4_source_44_source_sel <= 0;
      _stream_conv2d_4_source_44_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_44_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_44_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_44_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_44_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_44_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_44_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_44_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_44_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_44_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_44_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_44_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_44_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_44_pat_stride_buf_3 <= 0;
      __variable_wdata_1343 <= 0;
      _stream_conv2d_4_source_44_source_ram_raddr <= 0;
      _stream_conv2d_4_source_45_source_mode <= 5'b0;
      _stream_conv2d_4_source_45_source_offset <= 0;
      _source_stream_conv2d_4_source_45_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_45_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_45_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_45_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_3 <= 0;
      _stream_conv2d_4_source_45_source_sel <= 0;
      _stream_conv2d_4_source_45_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_45_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_45_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_45_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_45_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_45_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_45_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_45_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_45_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_45_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_45_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_45_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_45_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_45_pat_stride_buf_3 <= 0;
      __variable_wdata_1344 <= 0;
      _stream_conv2d_4_source_45_source_ram_raddr <= 0;
      _stream_conv2d_4_source_46_source_mode <= 5'b0;
      _stream_conv2d_4_source_46_source_offset <= 0;
      _source_stream_conv2d_4_source_46_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_46_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_46_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_46_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_3 <= 0;
      _stream_conv2d_4_source_46_source_sel <= 0;
      _stream_conv2d_4_source_46_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_46_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_46_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_46_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_46_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_46_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_46_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_46_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_46_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_46_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_46_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_46_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_46_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_46_pat_stride_buf_3 <= 0;
      __variable_wdata_1345 <= 0;
      _stream_conv2d_4_source_46_source_ram_raddr <= 0;
      _tmp_377 <= 0;
      _tmp_378 <= 0;
      _tmp_379 <= 0;
      _tmp_380 <= 0;
      _tmp_381 <= 0;
      _tmp_382 <= 0;
      _tmp_383 <= 0;
      _tmp_384 <= 0;
      _tmp_385 <= 0;
      _tmp_386 <= 0;
      _tmp_387 <= 0;
      _tmp_388 <= 0;
      _tmp_389 <= 0;
      _tmp_390 <= 0;
      _tmp_391 <= 0;
      _tmp_392 <= 0;
      _tmp_393 <= 0;
      _tmp_394 <= 0;
      _tmp_395 <= 0;
      _tmp_396 <= 0;
      _tmp_397 <= 0;
      _tmp_398 <= 0;
      _tmp_399 <= 0;
      _tmp_400 <= 0;
      _tmp_401 <= 0;
      _tmp_402 <= 0;
      _tmp_403 <= 0;
      _tmp_404 <= 0;
      _tmp_405 <= 0;
      _tmp_406 <= 0;
      _tmp_407 <= 0;
      _tmp_408 <= 0;
      _tmp_409 <= 0;
      _tmp_410 <= 0;
      _tmp_411 <= 0;
      _tmp_412 <= 0;
      _tmp_415 <= 0;
      _tmp_416 <= 0;
      _tmp_417 <= 0;
      _tmp_418 <= 0;
      _tmp_419 <= 0;
      _tmp_420 <= 0;
      _tmp_421 <= 0;
      _tmp_422 <= 0;
      _tmp_423 <= 0;
      _tmp_424 <= 0;
      _tmp_425 <= 0;
      _tmp_426 <= 0;
      _tmp_427 <= 0;
      _tmp_428 <= 0;
      _tmp_429 <= 0;
      _tmp_430 <= 0;
      _tmp_431 <= 0;
      _tmp_432 <= 0;
      _tmp_433 <= 0;
      _tmp_434 <= 0;
      _tmp_435 <= 0;
      _tmp_436 <= 0;
      _tmp_437 <= 0;
      _tmp_438 <= 0;
      _tmp_439 <= 0;
      _tmp_440 <= 0;
      _tmp_441 <= 0;
      _tmp_442 <= 0;
      _tmp_443 <= 0;
      _tmp_444 <= 0;
      _tmp_445 <= 0;
      _tmp_446 <= 0;
      _tmp_447 <= 0;
      _tmp_448 <= 0;
      _tmp_449 <= 0;
      _tmp_450 <= 0;
      _tmp_451 <= 0;
      _tmp_452 <= 0;
      _tmp_453 <= 0;
      _tmp_454 <= 0;
      _tmp_455 <= 0;
      _tmp_456 <= 0;
      _tmp_457 <= 0;
      _tmp_458 <= 0;
      _tmp_459 <= 0;
      _tmp_460 <= 0;
      _tmp_461 <= 0;
      _tmp_462 <= 0;
      _tmp_463 <= 0;
      _tmp_464 <= 0;
      _tmp_465 <= 0;
      _tmp_466 <= 0;
      _tmp_467 <= 0;
      _tmp_468 <= 0;
      _tmp_469 <= 0;
      _tmp_470 <= 0;
      _tmp_471 <= 0;
      _tmp_472 <= 0;
      _tmp_473 <= 0;
      _tmp_474 <= 0;
      _tmp_475 <= 0;
      _tmp_476 <= 0;
      _tmp_477 <= 0;
      _tmp_478 <= 0;
      _tmp_479 <= 0;
      _tmp_480 <= 0;
      _tmp_481 <= 0;
      _tmp_482 <= 0;
      _tmp_483 <= 0;
      _tmp_484 <= 0;
      _tmp_485 <= 0;
      _tmp_486 <= 0;
      _stream_conv2d_4_sink_89_sink_mode <= 5'b0;
      _stream_conv2d_4_sink_89_sink_offset <= 0;
      _stream_conv2d_4_sink_89_sink_size <= 0;
      _stream_conv2d_4_sink_89_sink_stride <= 0;
      _stream_conv2d_4_sink_89_sink_sel <= 0;
      _stream_conv2d_4_sink_89_sink_offset_buf <= 0;
      _stream_conv2d_4_sink_89_sink_size_buf <= 0;
      _stream_conv2d_4_sink_89_sink_stride_buf <= 0;
      _stream_conv2d_4_sink_89_sink_waddr <= 0;
      _stream_conv2d_4_sink_89_sink_count <= 0;
      _stream_conv2d_4_sink_89_sink_wdata <= 0;
      _tmp_1882 <= 0;
      _tmp_1883 <= 0;
      _tmp_1884 <= 0;
      _tmp_1885 <= 0;
      _tmp_1886 <= 0;
      _tmp_1887 <= 0;
      __variable_wdata_951 <= 0;
      _tmp_1888 <= 0;
      _tmp_1889 <= 0;
      _tmp_1890 <= 0;
      _tmp_1891 <= 0;
      _tmp_1894 <= 0;
      _tmp_1897 <= 0;
      _tmp_1898 <= 0;
      _tmp_1899 <= 0;
      _tmp_1900 <= 0;
      _tmp_1901 <= 0;
      _tmp_1902 <= 0;
      _tmp_1903 <= 0;
      _tmp_1904 <= 0;
      _tmp_1905 <= 0;
      _tmp_1906 <= 0;
      _tmp_1907 <= 0;
      _tmp_1908 <= 0;
      _tmp_1909 <= 0;
      _tmp_1910 <= 0;
      _tmp_1911 <= 0;
      _tmp_1912 <= 0;
      _tmp_1913 <= 0;
      _tmp_1914 <= 0;
      _tmp_1915 <= 0;
      _tmp_1916 <= 0;
      _tmp_1917 <= 0;
      _tmp_1918 <= 0;
      _tmp_1919 <= 0;
      _tmp_1920 <= 0;
      _tmp_1921 <= 0;
      _tmp_1922 <= 0;
      _tmp_1923 <= 0;
      _tmp_1924 <= 0;
      _tmp_1925 <= 0;
      _tmp_1926 <= 0;
      _tmp_1927 <= 0;
      _tmp_1928 <= 0;
      _tmp_1929 <= 0;
      _tmp_1930 <= 0;
      _tmp_1931 <= 0;
      _tmp_1932 <= 0;
      _tmp_1933 <= 0;
      _tmp_1934 <= 0;
      _tmp_1935 <= 0;
      _tmp_1936 <= 0;
      _tmp_1937 <= 0;
      _tmp_1938 <= 0;
      _tmp_1939 <= 0;
      _tmp_1940 <= 0;
      _tmp_1941 <= 0;
      _tmp_1942 <= 0;
      _tmp_1943 <= 0;
      _tmp_1944 <= 0;
      _tmp_1945 <= 0;
      _tmp_1946 <= 0;
      _tmp_1947 <= 0;
      _tmp_1948 <= 0;
      _tmp_1949 <= 0;
      _tmp_1950 <= 0;
      _tmp_1951 <= 0;
      _tmp_1952 <= 0;
      _tmp_1953 <= 0;
      _tmp_1954 <= 0;
      _tmp_1955 <= 0;
      _tmp_1956 <= 0;
      _tmp_1957 <= 0;
      _tmp_1958 <= 0;
      _tmp_1959 <= 0;
      _tmp_1960 <= 0;
      _tmp_1961 <= 0;
      _tmp_1962 <= 0;
      _tmp_1963 <= 0;
      _tmp_1964 <= 0;
      _tmp_1965 <= 0;
      _tmp_1966 <= 0;
      _tmp_1967 <= 0;
      _tmp_1968 <= 0;
      _tmp_1969 <= 0;
      _tmp_1970 <= 0;
      _tmp_1971 <= 0;
      _tmp_1972 <= 0;
      _tmp_1973 <= 0;
      _tmp_1974 <= 0;
      _tmp_1975 <= 0;
      _tmp_1976 <= 0;
      _tmp_1977 <= 0;
      _tmp_1978 <= 0;
      _tmp_1979 <= 0;
      _tmp_1980 <= 0;
      _tmp_1981 <= 0;
      _tmp_1982 <= 0;
      _tmp_1983 <= 0;
      _tmp_1984 <= 0;
      _tmp_1985 <= 0;
      _tmp_1986 <= 0;
      _tmp_1987 <= 0;
      _tmp_1988 <= 0;
      _tmp_1989 <= 0;
      _tmp_1990 <= 0;
      _tmp_1991 <= 0;
      _tmp_1992 <= 0;
      _tmp_1993 <= 0;
      _tmp_1994 <= 0;
      _tmp_1995 <= 0;
      _tmp_1996 <= 0;
      _tmp_1997 <= 0;
      _tmp_1998 <= 0;
      _tmp_1999 <= 0;
      _tmp_2000 <= 0;
      _tmp_2001 <= 0;
      _tmp_2002 <= 0;
      _tmp_2003 <= 0;
      _tmp_2004 <= 0;
      _tmp_2005 <= 0;
      _tmp_2006 <= 0;
      _stream_conv2d_4_busy_reg <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_7_idle <= _stream_conv2d_4_source_7_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_9_idle <= _stream_conv2d_4_source_9_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_11_source_ram_renable <= 0;
        _stream_conv2d_4_source_11_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_11_idle <= _stream_conv2d_4_source_11_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_13_source_ram_renable <= 0;
        _stream_conv2d_4_source_13_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_13_idle <= _stream_conv2d_4_source_13_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_15_source_ram_renable <= 0;
        _stream_conv2d_4_source_15_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_15_idle <= _stream_conv2d_4_source_15_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_20_idle <= _stream_conv2d_4_source_20_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_21_idle <= _stream_conv2d_4_source_21_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_22_idle <= _stream_conv2d_4_source_22_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_23_idle <= _stream_conv2d_4_source_23_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_24_idle <= _stream_conv2d_4_source_24_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_25_idle <= _stream_conv2d_4_source_25_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_26_idle <= _stream_conv2d_4_source_26_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_27_idle <= _stream_conv2d_4_source_27_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_28_idle <= _stream_conv2d_4_source_28_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_29_idle <= _stream_conv2d_4_source_29_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_30_idle <= _stream_conv2d_4_source_30_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_31_idle <= _stream_conv2d_4_source_31_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_32_idle <= _stream_conv2d_4_source_32_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_33_idle <= _stream_conv2d_4_source_33_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_34_idle <= _stream_conv2d_4_source_34_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_35_idle <= _stream_conv2d_4_source_35_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_36_idle <= _stream_conv2d_4_source_36_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_37_idle <= _stream_conv2d_4_source_37_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_38_source_ram_renable <= 0;
        _stream_conv2d_4_source_38_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_38_idle <= _stream_conv2d_4_source_38_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_39_source_ram_renable <= 0;
        _stream_conv2d_4_source_39_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_39_idle <= _stream_conv2d_4_source_39_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_40_source_ram_renable <= 0;
        _stream_conv2d_4_source_40_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_40_idle <= _stream_conv2d_4_source_40_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_41_source_ram_renable <= 0;
        _stream_conv2d_4_source_41_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_41_idle <= _stream_conv2d_4_source_41_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_42_source_ram_renable <= 0;
        _stream_conv2d_4_source_42_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_42_idle <= _stream_conv2d_4_source_42_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_43_source_ram_renable <= 0;
        _stream_conv2d_4_source_43_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_43_idle <= _stream_conv2d_4_source_43_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_44_source_ram_renable <= 0;
        _stream_conv2d_4_source_44_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_44_idle <= _stream_conv2d_4_source_44_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_45_source_ram_renable <= 0;
        _stream_conv2d_4_source_45_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_45_idle <= _stream_conv2d_4_source_45_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_46_source_ram_renable <= 0;
        _stream_conv2d_4_source_46_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_46_idle <= _stream_conv2d_4_source_46_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_89_sink_wenable <= 0;
        _stream_conv2d_4_sink_89_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_90_sink_wenable <= 0;
        _stream_conv2d_4_sink_90_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_1 <= _stream_conv2d_4_stream_ivalid;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_2 <= __stream_conv2d_4_stream_ivalid_1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_3 <= __stream_conv2d_4_stream_ivalid_2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_4 <= __stream_conv2d_4_stream_ivalid_3;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_5 <= __stream_conv2d_4_stream_ivalid_4;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_6 <= __stream_conv2d_4_stream_ivalid_5;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_7 <= __stream_conv2d_4_stream_ivalid_6;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_8 <= __stream_conv2d_4_stream_ivalid_7;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_9 <= __stream_conv2d_4_stream_ivalid_8;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_10 <= __stream_conv2d_4_stream_ivalid_9;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_11 <= __stream_conv2d_4_stream_ivalid_10;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_12 <= __stream_conv2d_4_stream_ivalid_11;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_13 <= __stream_conv2d_4_stream_ivalid_12;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_14 <= __stream_conv2d_4_stream_ivalid_13;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_15 <= __stream_conv2d_4_stream_ivalid_14;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_16 <= __stream_conv2d_4_stream_ivalid_15;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_17 <= __stream_conv2d_4_stream_ivalid_16;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_18 <= __stream_conv2d_4_stream_ivalid_17;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_19 <= __stream_conv2d_4_stream_ivalid_18;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_20 <= __stream_conv2d_4_stream_ivalid_19;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_21 <= __stream_conv2d_4_stream_ivalid_20;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_22 <= __stream_conv2d_4_stream_ivalid_21;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_23 <= __stream_conv2d_4_stream_ivalid_22;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_24 <= __stream_conv2d_4_stream_ivalid_23;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_25 <= __stream_conv2d_4_stream_ivalid_24;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_26 <= __stream_conv2d_4_stream_ivalid_25;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_27 <= __stream_conv2d_4_stream_ivalid_26;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_28 <= __stream_conv2d_4_stream_ivalid_27;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_29 <= __stream_conv2d_4_stream_ivalid_28;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_30 <= __stream_conv2d_4_stream_ivalid_29;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_31 <= __stream_conv2d_4_stream_ivalid_30;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_32 <= __stream_conv2d_4_stream_ivalid_31;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_33 <= __stream_conv2d_4_stream_ivalid_32;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_34 <= __stream_conv2d_4_stream_ivalid_33;
      end 
      if(_stream_conv2d_4_stream_ivalid && _stream_conv2d_4_stream_oready && _counter_reset_cond_952) begin
        _counter_data_952 <= 1'sd0;
      end 
      if(_stream_conv2d_4_stream_ivalid && _stream_conv2d_4_stream_oready) begin
        _counter_data_952 <= _counter_current_count_952;
      end 
      if(_stream_conv2d_4_stream_ivalid && _stream_conv2d_4_stream_oready) begin
        _counter_count_952 <= (_counter_current_count_952 >= stream_conv2d_4_parameter_0_data - 2'sd1)? _counter_current_count_952 + 2'sd1 - stream_conv2d_4_parameter_0_data : _counter_current_count_952 + 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _minus_data_957 <= stream_conv2d_4_parameter_0_data - 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _minus_data_963 <= stream_conv2d_4_parameter_0_data - 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1040 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1044 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1047 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1050 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1054 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1057 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1060 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1064 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1067 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1070 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1074 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1077 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1080 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1084 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1087 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1090 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1094 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1097 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1100 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1104 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1107 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1110 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1114 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1117 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1120 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1124 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1127 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1130 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1134 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1137 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1140 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1144 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1147 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1150 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1154 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1157 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1160 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1164 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1167 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1170 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1174 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1177 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1180 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1184 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1187 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1190 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1194 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1197 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1200 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1204 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1207 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1210 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1214 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1217 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1615 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1634 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1653 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1672 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1691 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1710 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1729 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1748 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1767 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1804 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1823 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1842 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1861 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1880 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1899 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1918 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1937 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1956 <= _cond_data_1001 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1972 <= _cond_data_1013 + stream_conv2d_4_parameter_17_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1991 <= _cond_data_1025 + stream_conv2d_4_parameter_18_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2033 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2052 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2071 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2090 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2109 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2128 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2147 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2166 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2185 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2222 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2241 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2260 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2279 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2298 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2317 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2336 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2355 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2374 <= _cond_data_1002 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2390 <= _cond_data_1014 + stream_conv2d_4_parameter_17_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2409 <= _cond_data_1026 + stream_conv2d_4_parameter_18_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2642_pointer_955 <= _pointer_data_955;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2644__variable_1033 <= stream_conv2d_4_source_22_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2645__variable_1032 <= stream_conv2d_4_source_21_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2646__variable_1031 <= stream_conv2d_4_source_20_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2647__variable_1036 <= stream_conv2d_4_source_25_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2648__variable_1035 <= stream_conv2d_4_source_24_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2649__variable_1034 <= stream_conv2d_4_source_23_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2650__variable_1039 <= stream_conv2d_4_source_28_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2651__variable_1038 <= stream_conv2d_4_source_27_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2652__variable_1037 <= stream_conv2d_4_source_26_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2655_pointer_1562 <= _pointer_data_1562;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2658_reinterpretcast_1349 <= _reinterpretcast_data_1349;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2663_pointer_961 <= _pointer_data_961;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2667_reinterpretcast_1353 <= _reinterpretcast_data_1353;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2674_pointer_1564 <= _pointer_data_1564;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2677_reinterpretcast_1357 <= _reinterpretcast_data_1357;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2684_reinterpretcast_1361 <= _reinterpretcast_data_1361;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2691_pointer_1566 <= _pointer_data_1566;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2694_reinterpretcast_1365 <= _reinterpretcast_data_1365;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2701_reinterpretcast_1369 <= _reinterpretcast_data_1369;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2708_pointer_1568 <= _pointer_data_1568;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2711_reinterpretcast_1373 <= _reinterpretcast_data_1373;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2718_reinterpretcast_1377 <= _reinterpretcast_data_1377;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2725_pointer_1570 <= _pointer_data_1570;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2728_reinterpretcast_1381 <= _reinterpretcast_data_1381;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2735_reinterpretcast_1385 <= _reinterpretcast_data_1385;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2742_pointer_1572 <= _pointer_data_1572;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2745_reinterpretcast_1389 <= _reinterpretcast_data_1389;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2752_reinterpretcast_1393 <= _reinterpretcast_data_1393;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2759_pointer_1574 <= _pointer_data_1574;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2762_reinterpretcast_1397 <= _reinterpretcast_data_1397;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2769_reinterpretcast_1401 <= _reinterpretcast_data_1401;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2776_pointer_1576 <= _pointer_data_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2779_reinterpretcast_1405 <= _reinterpretcast_data_1405;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2786_reinterpretcast_1409 <= _reinterpretcast_data_1409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2793_pointer_1578 <= _pointer_data_1578;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2796_reinterpretcast_1413 <= _reinterpretcast_data_1413;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2803_reinterpretcast_1417 <= _reinterpretcast_data_1417;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2808__variable_951 <= stream_conv2d_4__reduce_reset_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2839__variable_946 <= stream_conv2d_4_parameter_0_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2855_reinterpretcast_1457 <= _reinterpretcast_data_1457;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2860_reinterpretcast_1461 <= _reinterpretcast_data_1461;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2865_reinterpretcast_1465 <= _reinterpretcast_data_1465;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2870_reinterpretcast_1469 <= _reinterpretcast_data_1469;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2875_reinterpretcast_1473 <= _reinterpretcast_data_1473;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2880_reinterpretcast_1477 <= _reinterpretcast_data_1477;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2885_reinterpretcast_1481 <= _reinterpretcast_data_1481;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2890_reinterpretcast_1485 <= _reinterpretcast_data_1485;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2895_reinterpretcast_1489 <= _reinterpretcast_data_1489;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2900_reinterpretcast_1493 <= _reinterpretcast_data_1493;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2905_reinterpretcast_1497 <= _reinterpretcast_data_1497;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2910_reinterpretcast_1501 <= _reinterpretcast_data_1501;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2915_reinterpretcast_1505 <= _reinterpretcast_data_1505;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2920_reinterpretcast_1509 <= _reinterpretcast_data_1509;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2925_reinterpretcast_1513 <= _reinterpretcast_data_1513;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2930_reinterpretcast_1517 <= _reinterpretcast_data_1517;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2935_reinterpretcast_1521 <= _reinterpretcast_data_1521;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2940_reinterpretcast_1525 <= _reinterpretcast_data_1525;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2960_cond_978 <= _cond_data_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2982_cond_990 <= _cond_data_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3028_cond_977 <= _cond_data_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3050_cond_989 <= _cond_data_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_959 <= _counter_data_952 == _minus_data_957;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_965 <= _counter_data_952 == _minus_data_963;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2643__delay_2642_pointer_955 <= __delay_data_2642_pointer_955;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2653_reinterpretcast_1223 <= _reinterpretcast_data_1223;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2656__delay_2655_pointer_1562 <= __delay_data_2655_pointer_1562;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2659__delay_2658_reinterpretcast_1349 <= __delay_data_2658_reinterpretcast_1349;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2661_plus_1615 <= _plus_data_1615;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2664__delay_2663_pointer_961 <= __delay_data_2663_pointer_961;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2665_reinterpretcast_1227 <= _reinterpretcast_data_1227;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2668__delay_2667_reinterpretcast_1353 <= __delay_data_2667_reinterpretcast_1353;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2670_plus_1804 <= _plus_data_1804;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2672_reinterpretcast_1231 <= _reinterpretcast_data_1231;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2675__delay_2674_pointer_1564 <= __delay_data_2674_pointer_1564;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2678__delay_2677_reinterpretcast_1357 <= __delay_data_2677_reinterpretcast_1357;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2680_plus_1634 <= _plus_data_1634;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2682_reinterpretcast_1235 <= _reinterpretcast_data_1235;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2685__delay_2684_reinterpretcast_1361 <= __delay_data_2684_reinterpretcast_1361;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2687_plus_1823 <= _plus_data_1823;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2689_reinterpretcast_1239 <= _reinterpretcast_data_1239;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2692__delay_2691_pointer_1566 <= __delay_data_2691_pointer_1566;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2695__delay_2694_reinterpretcast_1365 <= __delay_data_2694_reinterpretcast_1365;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2697_plus_1653 <= _plus_data_1653;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2699_reinterpretcast_1243 <= _reinterpretcast_data_1243;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2702__delay_2701_reinterpretcast_1369 <= __delay_data_2701_reinterpretcast_1369;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2704_plus_1842 <= _plus_data_1842;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2706_reinterpretcast_1247 <= _reinterpretcast_data_1247;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2709__delay_2708_pointer_1568 <= __delay_data_2708_pointer_1568;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2712__delay_2711_reinterpretcast_1373 <= __delay_data_2711_reinterpretcast_1373;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2714_plus_1672 <= _plus_data_1672;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2716_reinterpretcast_1251 <= _reinterpretcast_data_1251;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2719__delay_2718_reinterpretcast_1377 <= __delay_data_2718_reinterpretcast_1377;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2721_plus_1861 <= _plus_data_1861;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2723_reinterpretcast_1255 <= _reinterpretcast_data_1255;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2726__delay_2725_pointer_1570 <= __delay_data_2725_pointer_1570;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2729__delay_2728_reinterpretcast_1381 <= __delay_data_2728_reinterpretcast_1381;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2731_plus_1691 <= _plus_data_1691;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2733_reinterpretcast_1259 <= _reinterpretcast_data_1259;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2736__delay_2735_reinterpretcast_1385 <= __delay_data_2735_reinterpretcast_1385;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2738_plus_1880 <= _plus_data_1880;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2740_reinterpretcast_1263 <= _reinterpretcast_data_1263;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2743__delay_2742_pointer_1572 <= __delay_data_2742_pointer_1572;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2746__delay_2745_reinterpretcast_1389 <= __delay_data_2745_reinterpretcast_1389;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2748_plus_1710 <= _plus_data_1710;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2750_reinterpretcast_1267 <= _reinterpretcast_data_1267;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2753__delay_2752_reinterpretcast_1393 <= __delay_data_2752_reinterpretcast_1393;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2755_plus_1899 <= _plus_data_1899;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2757_reinterpretcast_1271 <= _reinterpretcast_data_1271;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2760__delay_2759_pointer_1574 <= __delay_data_2759_pointer_1574;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2763__delay_2762_reinterpretcast_1397 <= __delay_data_2762_reinterpretcast_1397;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2765_plus_1729 <= _plus_data_1729;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2767_reinterpretcast_1275 <= _reinterpretcast_data_1275;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2770__delay_2769_reinterpretcast_1401 <= __delay_data_2769_reinterpretcast_1401;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2772_plus_1918 <= _plus_data_1918;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2774_reinterpretcast_1279 <= _reinterpretcast_data_1279;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2777__delay_2776_pointer_1576 <= __delay_data_2776_pointer_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2780__delay_2779_reinterpretcast_1405 <= __delay_data_2779_reinterpretcast_1405;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2782_plus_1748 <= _plus_data_1748;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2784_reinterpretcast_1283 <= _reinterpretcast_data_1283;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2787__delay_2786_reinterpretcast_1409 <= __delay_data_2786_reinterpretcast_1409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2789_plus_1937 <= _plus_data_1937;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2791_reinterpretcast_1287 <= _reinterpretcast_data_1287;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2794__delay_2793_pointer_1578 <= __delay_data_2793_pointer_1578;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2797__delay_2796_reinterpretcast_1413 <= __delay_data_2796_reinterpretcast_1413;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2799_plus_1767 <= _plus_data_1767;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2801_reinterpretcast_1291 <= _reinterpretcast_data_1291;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2804__delay_2803_reinterpretcast_1417 <= __delay_data_2803_reinterpretcast_1417;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2806_plus_1956 <= _plus_data_1956;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2809__delay_2808__variable_951 <= __delay_data_2808__variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2824_plus_1972 <= _plus_data_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2840__delay_2839__variable_946 <= __delay_data_2839__variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2856__delay_2855_reinterpretcast_1457 <= __delay_data_2855_reinterpretcast_1457;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2858_plus_2033 <= _plus_data_2033;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2861__delay_2860_reinterpretcast_1461 <= __delay_data_2860_reinterpretcast_1461;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2863_plus_2222 <= _plus_data_2222;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2866__delay_2865_reinterpretcast_1465 <= __delay_data_2865_reinterpretcast_1465;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2868_plus_2052 <= _plus_data_2052;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2871__delay_2870_reinterpretcast_1469 <= __delay_data_2870_reinterpretcast_1469;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2873_plus_2241 <= _plus_data_2241;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2876__delay_2875_reinterpretcast_1473 <= __delay_data_2875_reinterpretcast_1473;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2878_plus_2071 <= _plus_data_2071;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2881__delay_2880_reinterpretcast_1477 <= __delay_data_2880_reinterpretcast_1477;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2883_plus_2260 <= _plus_data_2260;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2886__delay_2885_reinterpretcast_1481 <= __delay_data_2885_reinterpretcast_1481;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2888_plus_2090 <= _plus_data_2090;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2891__delay_2890_reinterpretcast_1485 <= __delay_data_2890_reinterpretcast_1485;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2893_plus_2279 <= _plus_data_2279;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2896__delay_2895_reinterpretcast_1489 <= __delay_data_2895_reinterpretcast_1489;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2898_plus_2109 <= _plus_data_2109;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2901__delay_2900_reinterpretcast_1493 <= __delay_data_2900_reinterpretcast_1493;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2903_plus_2298 <= _plus_data_2298;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2906__delay_2905_reinterpretcast_1497 <= __delay_data_2905_reinterpretcast_1497;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2908_plus_2128 <= _plus_data_2128;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2911__delay_2910_reinterpretcast_1501 <= __delay_data_2910_reinterpretcast_1501;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2913_plus_2317 <= _plus_data_2317;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2916__delay_2915_reinterpretcast_1505 <= __delay_data_2915_reinterpretcast_1505;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2918_plus_2147 <= _plus_data_2147;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2921__delay_2920_reinterpretcast_1509 <= __delay_data_2920_reinterpretcast_1509;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2923_plus_2336 <= _plus_data_2336;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2926__delay_2925_reinterpretcast_1513 <= __delay_data_2925_reinterpretcast_1513;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2928_plus_2166 <= _plus_data_2166;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2931__delay_2930_reinterpretcast_1517 <= __delay_data_2930_reinterpretcast_1517;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2933_plus_2355 <= _plus_data_2355;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2936__delay_2935_reinterpretcast_1521 <= __delay_data_2935_reinterpretcast_1521;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2938_plus_2185 <= _plus_data_2185;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2941__delay_2940_reinterpretcast_1525 <= __delay_data_2940_reinterpretcast_1525;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2943_plus_2374 <= _plus_data_2374;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2945_plus_2390 <= _plus_data_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2961__delay_2960_cond_978 <= __delay_data_2960_cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2983__delay_2982_cond_990 <= __delay_data_2982_cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3005_plus_2409 <= _plus_data_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3029__delay_3028_cond_977 <= __delay_data_3028_cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3051__delay_3050_cond_989 <= __delay_data_3050_cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3073_plus_1991 <= _plus_data_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _land_data_960 <= __delay_data_2643__delay_2642_pointer_955 && _eq_data_959;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _land_data_966 <= __delay_data_2664__delay_2663_pointer_961 && _eq_data_965;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2654__delay_2653_reinterpretcast_1223 <= __delay_data_2653_reinterpretcast_1223;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2657__delay_2656__delay_2655_pointer_1562 <= __delay_data_2656__delay_2655_pointer_1562;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2660__delay_2659__delay_2658_reinterpretcast_1349 <= __delay_data_2659__delay_2658_reinterpretcast_1349;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2662__delay_2661_plus_1615 <= __delay_data_2661_plus_1615;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2666__delay_2665_reinterpretcast_1227 <= __delay_data_2665_reinterpretcast_1227;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2669__delay_2668__delay_2667_reinterpretcast_1353 <= __delay_data_2668__delay_2667_reinterpretcast_1353;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2671__delay_2670_plus_1804 <= __delay_data_2670_plus_1804;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2673__delay_2672_reinterpretcast_1231 <= __delay_data_2672_reinterpretcast_1231;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2676__delay_2675__delay_2674_pointer_1564 <= __delay_data_2675__delay_2674_pointer_1564;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2679__delay_2678__delay_2677_reinterpretcast_1357 <= __delay_data_2678__delay_2677_reinterpretcast_1357;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2681__delay_2680_plus_1634 <= __delay_data_2680_plus_1634;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2683__delay_2682_reinterpretcast_1235 <= __delay_data_2682_reinterpretcast_1235;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2686__delay_2685__delay_2684_reinterpretcast_1361 <= __delay_data_2685__delay_2684_reinterpretcast_1361;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2688__delay_2687_plus_1823 <= __delay_data_2687_plus_1823;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2690__delay_2689_reinterpretcast_1239 <= __delay_data_2689_reinterpretcast_1239;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2693__delay_2692__delay_2691_pointer_1566 <= __delay_data_2692__delay_2691_pointer_1566;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2696__delay_2695__delay_2694_reinterpretcast_1365 <= __delay_data_2695__delay_2694_reinterpretcast_1365;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2698__delay_2697_plus_1653 <= __delay_data_2697_plus_1653;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2700__delay_2699_reinterpretcast_1243 <= __delay_data_2699_reinterpretcast_1243;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2703__delay_2702__delay_2701_reinterpretcast_1369 <= __delay_data_2702__delay_2701_reinterpretcast_1369;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2705__delay_2704_plus_1842 <= __delay_data_2704_plus_1842;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2707__delay_2706_reinterpretcast_1247 <= __delay_data_2706_reinterpretcast_1247;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2710__delay_2709__delay_2708_pointer_1568 <= __delay_data_2709__delay_2708_pointer_1568;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2713__delay_2712__delay_2711_reinterpretcast_1373 <= __delay_data_2712__delay_2711_reinterpretcast_1373;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2715__delay_2714_plus_1672 <= __delay_data_2714_plus_1672;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2717__delay_2716_reinterpretcast_1251 <= __delay_data_2716_reinterpretcast_1251;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2720__delay_2719__delay_2718_reinterpretcast_1377 <= __delay_data_2719__delay_2718_reinterpretcast_1377;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2722__delay_2721_plus_1861 <= __delay_data_2721_plus_1861;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2724__delay_2723_reinterpretcast_1255 <= __delay_data_2723_reinterpretcast_1255;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2727__delay_2726__delay_2725_pointer_1570 <= __delay_data_2726__delay_2725_pointer_1570;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2730__delay_2729__delay_2728_reinterpretcast_1381 <= __delay_data_2729__delay_2728_reinterpretcast_1381;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2732__delay_2731_plus_1691 <= __delay_data_2731_plus_1691;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2734__delay_2733_reinterpretcast_1259 <= __delay_data_2733_reinterpretcast_1259;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2737__delay_2736__delay_2735_reinterpretcast_1385 <= __delay_data_2736__delay_2735_reinterpretcast_1385;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2739__delay_2738_plus_1880 <= __delay_data_2738_plus_1880;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2741__delay_2740_reinterpretcast_1263 <= __delay_data_2740_reinterpretcast_1263;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2744__delay_2743__delay_2742_pointer_1572 <= __delay_data_2743__delay_2742_pointer_1572;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2747__delay_2746__delay_2745_reinterpretcast_1389 <= __delay_data_2746__delay_2745_reinterpretcast_1389;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2749__delay_2748_plus_1710 <= __delay_data_2748_plus_1710;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2751__delay_2750_reinterpretcast_1267 <= __delay_data_2750_reinterpretcast_1267;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2754__delay_2753__delay_2752_reinterpretcast_1393 <= __delay_data_2753__delay_2752_reinterpretcast_1393;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2756__delay_2755_plus_1899 <= __delay_data_2755_plus_1899;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2758__delay_2757_reinterpretcast_1271 <= __delay_data_2757_reinterpretcast_1271;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2761__delay_2760__delay_2759_pointer_1574 <= __delay_data_2760__delay_2759_pointer_1574;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2764__delay_2763__delay_2762_reinterpretcast_1397 <= __delay_data_2763__delay_2762_reinterpretcast_1397;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2766__delay_2765_plus_1729 <= __delay_data_2765_plus_1729;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2768__delay_2767_reinterpretcast_1275 <= __delay_data_2767_reinterpretcast_1275;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2771__delay_2770__delay_2769_reinterpretcast_1401 <= __delay_data_2770__delay_2769_reinterpretcast_1401;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2773__delay_2772_plus_1918 <= __delay_data_2772_plus_1918;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2775__delay_2774_reinterpretcast_1279 <= __delay_data_2774_reinterpretcast_1279;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2778__delay_2777__delay_2776_pointer_1576 <= __delay_data_2777__delay_2776_pointer_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2781__delay_2780__delay_2779_reinterpretcast_1405 <= __delay_data_2780__delay_2779_reinterpretcast_1405;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2783__delay_2782_plus_1748 <= __delay_data_2782_plus_1748;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2785__delay_2784_reinterpretcast_1283 <= __delay_data_2784_reinterpretcast_1283;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2788__delay_2787__delay_2786_reinterpretcast_1409 <= __delay_data_2787__delay_2786_reinterpretcast_1409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2790__delay_2789_plus_1937 <= __delay_data_2789_plus_1937;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2792__delay_2791_reinterpretcast_1287 <= __delay_data_2791_reinterpretcast_1287;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2795__delay_2794__delay_2793_pointer_1578 <= __delay_data_2794__delay_2793_pointer_1578;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2798__delay_2797__delay_2796_reinterpretcast_1413 <= __delay_data_2797__delay_2796_reinterpretcast_1413;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2800__delay_2799_plus_1767 <= __delay_data_2799_plus_1767;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2802__delay_2801_reinterpretcast_1291 <= __delay_data_2801_reinterpretcast_1291;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2805__delay_2804__delay_2803_reinterpretcast_1417 <= __delay_data_2804__delay_2803_reinterpretcast_1417;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2807__delay_2806_plus_1956 <= __delay_data_2806_plus_1956;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2810__delay_2809__delay_2808__variable_951 <= __delay_data_2809__delay_2808__variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2825__delay_2824_plus_1972 <= __delay_data_2824_plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2841__delay_2840__delay_2839__variable_946 <= __delay_data_2840__delay_2839__variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2857__delay_2856__delay_2855_reinterpretcast_1457 <= __delay_data_2856__delay_2855_reinterpretcast_1457;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2859__delay_2858_plus_2033 <= __delay_data_2858_plus_2033;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2862__delay_2861__delay_2860_reinterpretcast_1461 <= __delay_data_2861__delay_2860_reinterpretcast_1461;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2864__delay_2863_plus_2222 <= __delay_data_2863_plus_2222;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2867__delay_2866__delay_2865_reinterpretcast_1465 <= __delay_data_2866__delay_2865_reinterpretcast_1465;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2869__delay_2868_plus_2052 <= __delay_data_2868_plus_2052;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2872__delay_2871__delay_2870_reinterpretcast_1469 <= __delay_data_2871__delay_2870_reinterpretcast_1469;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2874__delay_2873_plus_2241 <= __delay_data_2873_plus_2241;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2877__delay_2876__delay_2875_reinterpretcast_1473 <= __delay_data_2876__delay_2875_reinterpretcast_1473;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2879__delay_2878_plus_2071 <= __delay_data_2878_plus_2071;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2882__delay_2881__delay_2880_reinterpretcast_1477 <= __delay_data_2881__delay_2880_reinterpretcast_1477;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2884__delay_2883_plus_2260 <= __delay_data_2883_plus_2260;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2887__delay_2886__delay_2885_reinterpretcast_1481 <= __delay_data_2886__delay_2885_reinterpretcast_1481;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2889__delay_2888_plus_2090 <= __delay_data_2888_plus_2090;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2892__delay_2891__delay_2890_reinterpretcast_1485 <= __delay_data_2891__delay_2890_reinterpretcast_1485;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2894__delay_2893_plus_2279 <= __delay_data_2893_plus_2279;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2897__delay_2896__delay_2895_reinterpretcast_1489 <= __delay_data_2896__delay_2895_reinterpretcast_1489;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2899__delay_2898_plus_2109 <= __delay_data_2898_plus_2109;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2902__delay_2901__delay_2900_reinterpretcast_1493 <= __delay_data_2901__delay_2900_reinterpretcast_1493;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2904__delay_2903_plus_2298 <= __delay_data_2903_plus_2298;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2907__delay_2906__delay_2905_reinterpretcast_1497 <= __delay_data_2906__delay_2905_reinterpretcast_1497;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2909__delay_2908_plus_2128 <= __delay_data_2908_plus_2128;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2912__delay_2911__delay_2910_reinterpretcast_1501 <= __delay_data_2911__delay_2910_reinterpretcast_1501;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2914__delay_2913_plus_2317 <= __delay_data_2913_plus_2317;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2917__delay_2916__delay_2915_reinterpretcast_1505 <= __delay_data_2916__delay_2915_reinterpretcast_1505;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2919__delay_2918_plus_2147 <= __delay_data_2918_plus_2147;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2922__delay_2921__delay_2920_reinterpretcast_1509 <= __delay_data_2921__delay_2920_reinterpretcast_1509;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2924__delay_2923_plus_2336 <= __delay_data_2923_plus_2336;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2927__delay_2926__delay_2925_reinterpretcast_1513 <= __delay_data_2926__delay_2925_reinterpretcast_1513;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2929__delay_2928_plus_2166 <= __delay_data_2928_plus_2166;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2932__delay_2931__delay_2930_reinterpretcast_1517 <= __delay_data_2931__delay_2930_reinterpretcast_1517;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2934__delay_2933_plus_2355 <= __delay_data_2933_plus_2355;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2937__delay_2936__delay_2935_reinterpretcast_1521 <= __delay_data_2936__delay_2935_reinterpretcast_1521;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2939__delay_2938_plus_2185 <= __delay_data_2938_plus_2185;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2942__delay_2941__delay_2940_reinterpretcast_1525 <= __delay_data_2941__delay_2940_reinterpretcast_1525;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2944__delay_2943_plus_2374 <= __delay_data_2943_plus_2374;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2946__delay_2945_plus_2390 <= __delay_data_2945_plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2962__delay_2961__delay_2960_cond_978 <= __delay_data_2961__delay_2960_cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2984__delay_2983__delay_2982_cond_990 <= __delay_data_2983__delay_2982_cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3006__delay_3005_plus_2409 <= __delay_data_3005_plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3030__delay_3029__delay_3028_cond_977 <= __delay_data_3029__delay_3028_cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3052__delay_3051__delay_3050_cond_989 <= __delay_data_3051__delay_3050_cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3074__delay_3073_plus_1991 <= __delay_data_3073_plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2811__delay_2810__delay_2809____variable_951 <= __delay_data_2810__delay_2809__delay_2808__variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2826__delay_2825__delay_2824_plus_1972 <= __delay_data_2825__delay_2824_plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2842__delay_2841__delay_2840____variable_946 <= __delay_data_2841__delay_2840__delay_2839__variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2947__delay_2946__delay_2945_plus_2390 <= __delay_data_2946__delay_2945_plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2963__delay_2962__delay_2961__delay_2960_cond_978 <= __delay_data_2962__delay_2961__delay_2960_cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2985__delay_2984__delay_2983__delay_2982_cond_990 <= __delay_data_2984__delay_2983__delay_2982_cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3007__delay_3006__delay_3005_plus_2409 <= __delay_data_3006__delay_3005_plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3031__delay_3030__delay_3029__delay_3028_cond_977 <= __delay_data_3030__delay_3029__delay_3028_cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3053__delay_3052__delay_3051__delay_3050_cond_989 <= __delay_data_3052__delay_3051__delay_3050_cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3075__delay_3074__delay_3073_plus_1991 <= __delay_data_3074__delay_3073_plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2812__delay_2811__delay_2810____variable_951 <= __delay_data_2811__delay_2810__delay_2809____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2827__delay_2826__delay_2825___plus_1972 <= __delay_data_2826__delay_2825__delay_2824_plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2843__delay_2842__delay_2841____variable_946 <= __delay_data_2842__delay_2841__delay_2840____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2948__delay_2947__delay_2946___plus_2390 <= __delay_data_2947__delay_2946__delay_2945_plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2964__delay_2963__delay_2962__delay_2961___cond_978 <= __delay_data_2963__delay_2962__delay_2961__delay_2960_cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2986__delay_2985__delay_2984__delay_2983___cond_990 <= __delay_data_2985__delay_2984__delay_2983__delay_2982_cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3008__delay_3007__delay_3006___plus_2409 <= __delay_data_3007__delay_3006__delay_3005_plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3032__delay_3031__delay_3030__delay_3029___cond_977 <= __delay_data_3031__delay_3030__delay_3029__delay_3028_cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3054__delay_3053__delay_3052__delay_3051___cond_989 <= __delay_data_3053__delay_3052__delay_3051__delay_3050_cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3076__delay_3075__delay_3074___plus_1991 <= __delay_data_3075__delay_3074__delay_3073_plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2813__delay_2812__delay_2811____variable_951 <= __delay_data_2812__delay_2811__delay_2810____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2828__delay_2827__delay_2826___plus_1972 <= __delay_data_2827__delay_2826__delay_2825___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2844__delay_2843__delay_2842____variable_946 <= __delay_data_2843__delay_2842__delay_2841____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2949__delay_2948__delay_2947___plus_2390 <= __delay_data_2948__delay_2947__delay_2946___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2965__delay_2964__delay_2963__delay_2962___cond_978 <= __delay_data_2964__delay_2963__delay_2962__delay_2961___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2987__delay_2986__delay_2985__delay_2984___cond_990 <= __delay_data_2986__delay_2985__delay_2984__delay_2983___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3009__delay_3008__delay_3007___plus_2409 <= __delay_data_3008__delay_3007__delay_3006___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3033__delay_3032__delay_3031__delay_3030___cond_977 <= __delay_data_3032__delay_3031__delay_3030__delay_3029___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3055__delay_3054__delay_3053__delay_3052___cond_989 <= __delay_data_3054__delay_3053__delay_3052__delay_3051___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3077__delay_3076__delay_3075___plus_1991 <= __delay_data_3076__delay_3075__delay_3074___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2814__delay_2813__delay_2812____variable_951 <= __delay_data_2813__delay_2812__delay_2811____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2829__delay_2828__delay_2827___plus_1972 <= __delay_data_2828__delay_2827__delay_2826___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2845__delay_2844__delay_2843____variable_946 <= __delay_data_2844__delay_2843__delay_2842____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2950__delay_2949__delay_2948___plus_2390 <= __delay_data_2949__delay_2948__delay_2947___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2966__delay_2965__delay_2964__delay_2963___cond_978 <= __delay_data_2965__delay_2964__delay_2963__delay_2962___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2988__delay_2987__delay_2986__delay_2985___cond_990 <= __delay_data_2987__delay_2986__delay_2985__delay_2984___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3010__delay_3009__delay_3008___plus_2409 <= __delay_data_3009__delay_3008__delay_3007___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3034__delay_3033__delay_3032__delay_3031___cond_977 <= __delay_data_3033__delay_3032__delay_3031__delay_3030___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3056__delay_3055__delay_3054__delay_3053___cond_989 <= __delay_data_3055__delay_3054__delay_3053__delay_3052___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3078__delay_3077__delay_3076___plus_1991 <= __delay_data_3077__delay_3076__delay_3075___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2815__delay_2814__delay_2813____variable_951 <= __delay_data_2814__delay_2813__delay_2812____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2830__delay_2829__delay_2828___plus_1972 <= __delay_data_2829__delay_2828__delay_2827___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2846__delay_2845__delay_2844____variable_946 <= __delay_data_2845__delay_2844__delay_2843____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2951__delay_2950__delay_2949___plus_2390 <= __delay_data_2950__delay_2949__delay_2948___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2967__delay_2966__delay_2965__delay_2964___cond_978 <= __delay_data_2966__delay_2965__delay_2964__delay_2963___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2989__delay_2988__delay_2987__delay_2986___cond_990 <= __delay_data_2988__delay_2987__delay_2986__delay_2985___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3011__delay_3010__delay_3009___plus_2409 <= __delay_data_3010__delay_3009__delay_3008___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3035__delay_3034__delay_3033__delay_3032___cond_977 <= __delay_data_3034__delay_3033__delay_3032__delay_3031___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3057__delay_3056__delay_3055__delay_3054___cond_989 <= __delay_data_3056__delay_3055__delay_3054__delay_3053___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3079__delay_3078__delay_3077___plus_1991 <= __delay_data_3078__delay_3077__delay_3076___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2816__delay_2815__delay_2814____variable_951 <= __delay_data_2815__delay_2814__delay_2813____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2831__delay_2830__delay_2829___plus_1972 <= __delay_data_2830__delay_2829__delay_2828___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2847__delay_2846__delay_2845____variable_946 <= __delay_data_2846__delay_2845__delay_2844____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2952__delay_2951__delay_2950___plus_2390 <= __delay_data_2951__delay_2950__delay_2949___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2968__delay_2967__delay_2966__delay_2965___cond_978 <= __delay_data_2967__delay_2966__delay_2965__delay_2964___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2990__delay_2989__delay_2988__delay_2987___cond_990 <= __delay_data_2989__delay_2988__delay_2987__delay_2986___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3012__delay_3011__delay_3010___plus_2409 <= __delay_data_3011__delay_3010__delay_3009___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3036__delay_3035__delay_3034__delay_3033___cond_977 <= __delay_data_3035__delay_3034__delay_3033__delay_3032___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3058__delay_3057__delay_3056__delay_3055___cond_989 <= __delay_data_3057__delay_3056__delay_3055__delay_3054___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3080__delay_3079__delay_3078___plus_1991 <= __delay_data_3079__delay_3078__delay_3077___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2817__delay_2816__delay_2815____variable_951 <= __delay_data_2816__delay_2815__delay_2814____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2832__delay_2831__delay_2830___plus_1972 <= __delay_data_2831__delay_2830__delay_2829___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2848__delay_2847__delay_2846____variable_946 <= __delay_data_2847__delay_2846__delay_2845____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2953__delay_2952__delay_2951___plus_2390 <= __delay_data_2952__delay_2951__delay_2950___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2969__delay_2968__delay_2967__delay_2966___cond_978 <= __delay_data_2968__delay_2967__delay_2966__delay_2965___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2991__delay_2990__delay_2989__delay_2988___cond_990 <= __delay_data_2990__delay_2989__delay_2988__delay_2987___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3013__delay_3012__delay_3011___plus_2409 <= __delay_data_3012__delay_3011__delay_3010___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3037__delay_3036__delay_3035__delay_3034___cond_977 <= __delay_data_3036__delay_3035__delay_3034__delay_3033___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3059__delay_3058__delay_3057__delay_3056___cond_989 <= __delay_data_3058__delay_3057__delay_3056__delay_3055___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3081__delay_3080__delay_3079___plus_1991 <= __delay_data_3080__delay_3079__delay_3078___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2818__delay_2817__delay_2816____variable_951 <= __delay_data_2817__delay_2816__delay_2815____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2833__delay_2832__delay_2831___plus_1972 <= __delay_data_2832__delay_2831__delay_2830___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2849__delay_2848__delay_2847____variable_946 <= __delay_data_2848__delay_2847__delay_2846____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2954__delay_2953__delay_2952___plus_2390 <= __delay_data_2953__delay_2952__delay_2951___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2970__delay_2969__delay_2968__delay_2967___cond_978 <= __delay_data_2969__delay_2968__delay_2967__delay_2966___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2992__delay_2991__delay_2990__delay_2989___cond_990 <= __delay_data_2991__delay_2990__delay_2989__delay_2988___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3014__delay_3013__delay_3012___plus_2409 <= __delay_data_3013__delay_3012__delay_3011___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3038__delay_3037__delay_3036__delay_3035___cond_977 <= __delay_data_3037__delay_3036__delay_3035__delay_3034___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3060__delay_3059__delay_3058__delay_3057___cond_989 <= __delay_data_3059__delay_3058__delay_3057__delay_3056___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3082__delay_3081__delay_3080___plus_1991 <= __delay_data_3081__delay_3080__delay_3079___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2819__delay_2818__delay_2817____variable_951 <= __delay_data_2818__delay_2817__delay_2816____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2834__delay_2833__delay_2832___plus_1972 <= __delay_data_2833__delay_2832__delay_2831___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2850__delay_2849__delay_2848____variable_946 <= __delay_data_2849__delay_2848__delay_2847____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2955__delay_2954__delay_2953___plus_2390 <= __delay_data_2954__delay_2953__delay_2952___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2971__delay_2970__delay_2969__delay_2968___cond_978 <= __delay_data_2970__delay_2969__delay_2968__delay_2967___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2993__delay_2992__delay_2991__delay_2990___cond_990 <= __delay_data_2992__delay_2991__delay_2990__delay_2989___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3015__delay_3014__delay_3013___plus_2409 <= __delay_data_3014__delay_3013__delay_3012___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3039__delay_3038__delay_3037__delay_3036___cond_977 <= __delay_data_3038__delay_3037__delay_3036__delay_3035___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3061__delay_3060__delay_3059__delay_3058___cond_989 <= __delay_data_3060__delay_3059__delay_3058__delay_3057___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3083__delay_3082__delay_3081___plus_1991 <= __delay_data_3082__delay_3081__delay_3080___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2820__delay_2819__delay_2818____variable_951 <= __delay_data_2819__delay_2818__delay_2817____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2835__delay_2834__delay_2833___plus_1972 <= __delay_data_2834__delay_2833__delay_2832___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2851__delay_2850__delay_2849____variable_946 <= __delay_data_2850__delay_2849__delay_2848____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2956__delay_2955__delay_2954___plus_2390 <= __delay_data_2955__delay_2954__delay_2953___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2972__delay_2971__delay_2970__delay_2969___cond_978 <= __delay_data_2971__delay_2970__delay_2969__delay_2968___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2994__delay_2993__delay_2992__delay_2991___cond_990 <= __delay_data_2993__delay_2992__delay_2991__delay_2990___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3016__delay_3015__delay_3014___plus_2409 <= __delay_data_3015__delay_3014__delay_3013___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3040__delay_3039__delay_3038__delay_3037___cond_977 <= __delay_data_3039__delay_3038__delay_3037__delay_3036___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3062__delay_3061__delay_3060__delay_3059___cond_989 <= __delay_data_3061__delay_3060__delay_3059__delay_3058___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3084__delay_3083__delay_3082___plus_1991 <= __delay_data_3083__delay_3082__delay_3081___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2821__delay_2820__delay_2819____variable_951 <= __delay_data_2820__delay_2819__delay_2818____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2836__delay_2835__delay_2834___plus_1972 <= __delay_data_2835__delay_2834__delay_2833___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2852__delay_2851__delay_2850____variable_946 <= __delay_data_2851__delay_2850__delay_2849____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2957__delay_2956__delay_2955___plus_2390 <= __delay_data_2956__delay_2955__delay_2954___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2973__delay_2972__delay_2971__delay_2970___cond_978 <= __delay_data_2972__delay_2971__delay_2970__delay_2969___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2995__delay_2994__delay_2993__delay_2992___cond_990 <= __delay_data_2994__delay_2993__delay_2992__delay_2991___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3017__delay_3016__delay_3015___plus_2409 <= __delay_data_3016__delay_3015__delay_3014___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3041__delay_3040__delay_3039__delay_3038___cond_977 <= __delay_data_3040__delay_3039__delay_3038__delay_3037___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3063__delay_3062__delay_3061__delay_3060___cond_989 <= __delay_data_3062__delay_3061__delay_3060__delay_3059___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3085__delay_3084__delay_3083___plus_1991 <= __delay_data_3084__delay_3083__delay_3082___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2822__delay_2821__delay_2820____variable_951 <= __delay_data_2821__delay_2820__delay_2819____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2837__delay_2836__delay_2835___plus_1972 <= __delay_data_2836__delay_2835__delay_2834___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2853__delay_2852__delay_2851____variable_946 <= __delay_data_2852__delay_2851__delay_2850____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2958__delay_2957__delay_2956___plus_2390 <= __delay_data_2957__delay_2956__delay_2955___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2974__delay_2973__delay_2972__delay_2971___cond_978 <= __delay_data_2973__delay_2972__delay_2971__delay_2970___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2996__delay_2995__delay_2994__delay_2993___cond_990 <= __delay_data_2995__delay_2994__delay_2993__delay_2992___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3018__delay_3017__delay_3016___plus_2409 <= __delay_data_3017__delay_3016__delay_3015___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3042__delay_3041__delay_3040__delay_3039___cond_977 <= __delay_data_3041__delay_3040__delay_3039__delay_3038___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3064__delay_3063__delay_3062__delay_3061___cond_989 <= __delay_data_3063__delay_3062__delay_3061__delay_3060___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3086__delay_3085__delay_3084___plus_1991 <= __delay_data_3085__delay_3084__delay_3083___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2823__delay_2822__delay_2821____variable_951 <= __delay_data_2822__delay_2821__delay_2820____variable_951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2838__delay_2837__delay_2836___plus_1972 <= __delay_data_2837__delay_2836__delay_2835___plus_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2854__delay_2853__delay_2852____variable_946 <= __delay_data_2853__delay_2852__delay_2851____variable_946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2959__delay_2958__delay_2957___plus_2390 <= __delay_data_2958__delay_2957__delay_2956___plus_2390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2975__delay_2974__delay_2973__delay_2972___cond_978 <= __delay_data_2974__delay_2973__delay_2972__delay_2971___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2997__delay_2996__delay_2995__delay_2994___cond_990 <= __delay_data_2996__delay_2995__delay_2994__delay_2993___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3019__delay_3018__delay_3017___plus_2409 <= __delay_data_3018__delay_3017__delay_3016___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3043__delay_3042__delay_3041__delay_3040___cond_977 <= __delay_data_3042__delay_3041__delay_3040__delay_3039___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3065__delay_3064__delay_3063__delay_3062___cond_989 <= __delay_data_3064__delay_3063__delay_3062__delay_3061___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3087__delay_3086__delay_3085___plus_1991 <= __delay_data_3086__delay_3085__delay_3084___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2976__delay_2975__delay_2974__delay_2973___cond_978 <= __delay_data_2975__delay_2974__delay_2973__delay_2972___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2998__delay_2997__delay_2996__delay_2995___cond_990 <= __delay_data_2997__delay_2996__delay_2995__delay_2994___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3020__delay_3019__delay_3018___plus_2409 <= __delay_data_3019__delay_3018__delay_3017___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3044__delay_3043__delay_3042__delay_3041___cond_977 <= __delay_data_3043__delay_3042__delay_3041__delay_3040___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3066__delay_3065__delay_3064__delay_3063___cond_989 <= __delay_data_3065__delay_3064__delay_3063__delay_3062___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3088__delay_3087__delay_3086___plus_1991 <= __delay_data_3087__delay_3086__delay_3085___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2977__delay_2976__delay_2975__delay_2974___cond_978 <= __delay_data_2976__delay_2975__delay_2974__delay_2973___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2999__delay_2998__delay_2997__delay_2996___cond_990 <= __delay_data_2998__delay_2997__delay_2996__delay_2995___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3021__delay_3020__delay_3019___plus_2409 <= __delay_data_3020__delay_3019__delay_3018___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3045__delay_3044__delay_3043__delay_3042___cond_977 <= __delay_data_3044__delay_3043__delay_3042__delay_3041___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3067__delay_3066__delay_3065__delay_3064___cond_989 <= __delay_data_3066__delay_3065__delay_3064__delay_3063___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3089__delay_3088__delay_3087___plus_1991 <= __delay_data_3088__delay_3087__delay_3086___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2978__delay_2977__delay_2976__delay_2975___cond_978 <= __delay_data_2977__delay_2976__delay_2975__delay_2974___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3000__delay_2999__delay_2998__delay_2997___cond_990 <= __delay_data_2999__delay_2998__delay_2997__delay_2996___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3022__delay_3021__delay_3020___plus_2409 <= __delay_data_3021__delay_3020__delay_3019___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3046__delay_3045__delay_3044__delay_3043___cond_977 <= __delay_data_3045__delay_3044__delay_3043__delay_3042___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3068__delay_3067__delay_3066__delay_3065___cond_989 <= __delay_data_3067__delay_3066__delay_3065__delay_3064___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3090__delay_3089__delay_3088___plus_1991 <= __delay_data_3089__delay_3088__delay_3087___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2979__delay_2978__delay_2977__delay_2976___cond_978 <= __delay_data_2978__delay_2977__delay_2976__delay_2975___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3001__delay_3000__delay_2999__delay_2998___cond_990 <= __delay_data_3000__delay_2999__delay_2998__delay_2997___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3023__delay_3022__delay_3021___plus_2409 <= __delay_data_3022__delay_3021__delay_3020___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3047__delay_3046__delay_3045__delay_3044___cond_977 <= __delay_data_3046__delay_3045__delay_3044__delay_3043___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3069__delay_3068__delay_3067__delay_3066___cond_989 <= __delay_data_3068__delay_3067__delay_3066__delay_3065___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3091__delay_3090__delay_3089___plus_1991 <= __delay_data_3090__delay_3089__delay_3088___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2980__delay_2979__delay_2978__delay_2977___cond_978 <= __delay_data_2979__delay_2978__delay_2977__delay_2976___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3002__delay_3001__delay_3000__delay_2999___cond_990 <= __delay_data_3001__delay_3000__delay_2999__delay_2998___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3024__delay_3023__delay_3022___plus_2409 <= __delay_data_3023__delay_3022__delay_3021___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3048__delay_3047__delay_3046__delay_3045___cond_977 <= __delay_data_3047__delay_3046__delay_3045__delay_3044___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3070__delay_3069__delay_3068__delay_3067___cond_989 <= __delay_data_3069__delay_3068__delay_3067__delay_3066___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3092__delay_3091__delay_3090___plus_1991 <= __delay_data_3091__delay_3090__delay_3089___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2981__delay_2980__delay_2979__delay_2978___cond_978 <= __delay_data_2980__delay_2979__delay_2978__delay_2977___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3003__delay_3002__delay_3001__delay_3000___cond_990 <= __delay_data_3002__delay_3001__delay_3000__delay_2999___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3025__delay_3024__delay_3023___plus_2409 <= __delay_data_3024__delay_3023__delay_3022___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3049__delay_3048__delay_3047__delay_3046___cond_977 <= __delay_data_3048__delay_3047__delay_3046__delay_3045___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3071__delay_3070__delay_3069__delay_3068___cond_989 <= __delay_data_3070__delay_3069__delay_3068__delay_3067___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3093__delay_3092__delay_3091___plus_1991 <= __delay_data_3092__delay_3091__delay_3090___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1975 <= __substreamoutput_data_1973 + __delay_data_3049__delay_3048__delay_3047__delay_3046___cond_977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2393 <= __substreamoutput_data_2391 + __delay_data_2981__delay_2980__delay_2979__delay_2978___cond_978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3004__delay_3003__delay_3002__delay_3001___cond_990 <= __delay_data_3003__delay_3002__delay_3001__delay_3000___cond_990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3026__delay_3025__delay_3024___plus_2409 <= __delay_data_3025__delay_3024__delay_3023___plus_2409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3072__delay_3071__delay_3070__delay_3069___cond_989 <= __delay_data_3071__delay_3070__delay_3069__delay_3068___cond_989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3094__delay_3093__delay_3092___plus_1991 <= __delay_data_3093__delay_3092__delay_3091___plus_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3096__substreamoutput_1974 <= __substreamoutput_data_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3097__delay_3096__substreamoutput_1974 <= __delay_data_3096__substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3098__delay_3097____substreamoutput_1974 <= __delay_data_3097__delay_3096__substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3099__delay_3098____substreamoutput_1974 <= __delay_data_3098__delay_3097____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3100__delay_3099____substreamoutput_1974 <= __delay_data_3099__delay_3098____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3101__delay_3100____substreamoutput_1974 <= __delay_data_3100__delay_3099____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3102__delay_3101____substreamoutput_1974 <= __delay_data_3101__delay_3100____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3103__delay_3102____substreamoutput_1974 <= __delay_data_3102__delay_3101____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3104__delay_3103____substreamoutput_1974 <= __delay_data_3103__delay_3102____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3105__delay_3104____substreamoutput_1974 <= __delay_data_3104__delay_3103____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _greaterthan_data_1994 <= __substreamoutput_data_1992 > 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _greaterthan_data_2412 <= __substreamoutput_data_2410 > 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3027__substreamoutput_2410 <= __substreamoutput_data_2410;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3095__substreamoutput_1992 <= __substreamoutput_data_1992;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3106__delay_3105____substreamoutput_1974 <= __delay_data_3105__delay_3104____substreamoutput_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _cond_data_1996 <= (_greaterthan_data_1994)? __delay_data_3095__substreamoutput_1992 : 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _cond_data_2414 <= (_greaterthan_data_2412)? __delay_data_3027__substreamoutput_2410 : 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_3107__delay_3106____substreamoutput_1974 <= __delay_data_3106__delay_3105____substreamoutput_1974;
      end 
      if(_set_flag_272) begin
        _stream_conv2d_4_parameter_0_next_parameter_data <= cparam_conv2d_4_stream_reduce_size;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_946 <= _stream_conv2d_4_parameter_0_next_parameter_data;
      end 
      if(_set_flag_273) begin
        _stream_conv2d_4_parameter_1_next_parameter_data <= conv2d_4_col_select;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_947 <= _stream_conv2d_4_parameter_1_next_parameter_data;
      end 
      if(_set_flag_274) begin
        _stream_conv2d_4_parameter_2_next_parameter_data <= conv2d_4_row_select_buf;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_948 <= _stream_conv2d_4_parameter_2_next_parameter_data;
      end 
      if(_set_flag_275) begin
        _stream_conv2d_4_parameter_3_next_parameter_data <= conv2d_4_stream_pad_masks;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_949 <= _stream_conv2d_4_parameter_3_next_parameter_data;
      end 
      if(_set_flag_276) begin
        _stream_conv2d_4_parameter_4_next_parameter_data <= cparam_conv2d_4_stream_omit_mask;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_950 <= _stream_conv2d_4_parameter_4_next_parameter_data;
      end 
      if(_set_flag_277) begin
        _stream_conv2d_4_parameter_6_next_parameter_data <= cparam_conv2d_4_bias_scala;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_967 <= _stream_conv2d_4_parameter_6_next_parameter_data;
      end 
      if(_set_flag_278) begin
        _stream_conv2d_4_source_7_source_mode <= 5'b10;
        _stream_conv2d_4_source_7_source_offset <= (cparam_conv2d_4_bias_num == 1)? 0 : conv2d_4_och_count_buf;
      end 
      if(_set_flag_278) begin
        _source_stream_conv2d_4_source_7_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_278) begin
        _source_stream_conv2d_4_source_7_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_7_pat_stride_1 <= (cparam_conv2d_4_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_278) begin
        _source_stream_conv2d_4_source_7_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_278) begin
        _source_stream_conv2d_4_source_7_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_278) begin
        _stream_conv2d_4_source_7_source_sel <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_offset_buf <= _stream_conv2d_4_source_7_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_0 <= _source_stream_conv2d_4_source_7_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_1 <= _source_stream_conv2d_4_source_7_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_2 <= _source_stream_conv2d_4_source_7_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_3 <= _source_stream_conv2d_4_source_7_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_0 <= _source_stream_conv2d_4_source_7_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_1 <= _source_stream_conv2d_4_source_7_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_2 <= _source_stream_conv2d_4_source_7_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_3 <= _source_stream_conv2d_4_source_7_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_968 <= _stream_conv2d_4_source_7_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_idle <= 0;
        _stream_conv2d_4_source_7_source_ram_raddr <= _stream_conv2d_4_source_7_source_pat_all_offset;
        _stream_conv2d_4_source_7_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= _source_stream_conv2d_4_source_7_pat_cur_offset_0 + _source_stream_conv2d_4_source_7_pat_stride_buf_0;
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= _source_stream_conv2d_4_source_7_pat_cur_offset_1 + _source_stream_conv2d_4_source_7_pat_stride_buf_1;
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= _source_stream_conv2d_4_source_7_pat_cur_offset_2 + _source_stream_conv2d_4_source_7_pat_stride_buf_2;
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= _source_stream_conv2d_4_source_7_pat_cur_offset_3 + _source_stream_conv2d_4_source_7_pat_stride_buf_3;
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_7_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_idle <= 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_idle <= 1;
      end 
      if(_set_flag_281) begin
        _stream_conv2d_4_parameter_8_next_parameter_data <= cparam_conv2d_4_scale_scala;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_979 <= _stream_conv2d_4_parameter_8_next_parameter_data;
      end 
      if(_set_flag_282) begin
        _stream_conv2d_4_source_9_source_mode <= 5'b10;
        _stream_conv2d_4_source_9_source_offset <= (cparam_conv2d_4_scale_num == 1)? 0 : conv2d_4_och_count_buf;
      end 
      if(_set_flag_282) begin
        _source_stream_conv2d_4_source_9_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_282) begin
        _source_stream_conv2d_4_source_9_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_9_pat_stride_1 <= (cparam_conv2d_4_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_282) begin
        _source_stream_conv2d_4_source_9_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_282) begin
        _source_stream_conv2d_4_source_9_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_282) begin
        _stream_conv2d_4_source_9_source_sel <= 2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_offset_buf <= _stream_conv2d_4_source_9_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_0 <= _source_stream_conv2d_4_source_9_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_1 <= _source_stream_conv2d_4_source_9_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_2 <= _source_stream_conv2d_4_source_9_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_3 <= _source_stream_conv2d_4_source_9_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_0 <= _source_stream_conv2d_4_source_9_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_1 <= _source_stream_conv2d_4_source_9_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_2 <= _source_stream_conv2d_4_source_9_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_3 <= _source_stream_conv2d_4_source_9_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_980 <= _stream_conv2d_4_source_9_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_idle <= 0;
        _stream_conv2d_4_source_9_source_ram_raddr <= _stream_conv2d_4_source_9_source_pat_all_offset;
        _stream_conv2d_4_source_9_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= _source_stream_conv2d_4_source_9_pat_cur_offset_0 + _source_stream_conv2d_4_source_9_pat_stride_buf_0;
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= _source_stream_conv2d_4_source_9_pat_cur_offset_1 + _source_stream_conv2d_4_source_9_pat_stride_buf_1;
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= _source_stream_conv2d_4_source_9_pat_cur_offset_2 + _source_stream_conv2d_4_source_9_pat_stride_buf_2;
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= _source_stream_conv2d_4_source_9_pat_cur_offset_3 + _source_stream_conv2d_4_source_9_pat_stride_buf_3;
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_9_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_idle <= 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_idle <= 1;
      end 
      if(_set_flag_285) begin
        _stream_conv2d_4_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_991 <= _stream_conv2d_4_parameter_10_next_parameter_data;
      end 
      if(_set_flag_286) begin
        _stream_conv2d_4_source_11_source_mode <= 5'b0;
        _stream_conv2d_4_source_11_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_11_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_11_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_11_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_992 <= _stream_conv2d_4_source_11_source_empty_data;
      end 
      if(_set_flag_287) begin
        _stream_conv2d_4_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1003 <= _stream_conv2d_4_parameter_12_next_parameter_data;
      end 
      if(_set_flag_288) begin
        _stream_conv2d_4_source_13_source_mode <= 5'b0;
        _stream_conv2d_4_source_13_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_13_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_13_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_13_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_1004 <= _stream_conv2d_4_source_13_source_empty_data;
      end 
      if(_set_flag_289) begin
        _stream_conv2d_4_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1015 <= _stream_conv2d_4_parameter_14_next_parameter_data;
      end 
      if(_set_flag_290) begin
        _stream_conv2d_4_source_15_source_mode <= 5'b0;
        _stream_conv2d_4_source_15_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_15_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_15_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_15_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_1016 <= _stream_conv2d_4_source_15_source_empty_data;
      end 
      if(_set_flag_291) begin
        _stream_conv2d_4_parameter_16_next_parameter_data <= cparam_conv2d_4_cshamt_mul_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1027 <= _stream_conv2d_4_parameter_16_next_parameter_data;
      end 
      if(_set_flag_292) begin
        _stream_conv2d_4_parameter_17_next_parameter_data <= cparam_conv2d_4_cshamt_sum_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1028 <= _stream_conv2d_4_parameter_17_next_parameter_data;
      end 
      if(_set_flag_293) begin
        _stream_conv2d_4_parameter_18_next_parameter_data <= cparam_conv2d_4_cshamt_out_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1029 <= _stream_conv2d_4_parameter_18_next_parameter_data;
      end 
      if(_set_flag_294) begin
        _stream_conv2d_4_parameter_19_next_parameter_data <= cparam_conv2d_4_act_func_index;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1030 <= _stream_conv2d_4_parameter_19_next_parameter_data;
      end 
      if(_set_flag_295) begin
        _stream_conv2d_4_source_20_source_mode <= 5'b10;
        _stream_conv2d_4_source_20_source_offset <= conv2d_4_stream_act_local_0 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_295) begin
        _source_stream_conv2d_4_source_20_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_295) begin
        _source_stream_conv2d_4_source_20_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_295) begin
        _source_stream_conv2d_4_source_20_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_295) begin
        _source_stream_conv2d_4_source_20_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_295) begin
        _stream_conv2d_4_source_20_source_sel <= 3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_offset_buf <= _stream_conv2d_4_source_20_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_0 <= _source_stream_conv2d_4_source_20_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_1 <= _source_stream_conv2d_4_source_20_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_2 <= _source_stream_conv2d_4_source_20_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_3 <= _source_stream_conv2d_4_source_20_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_0 <= _source_stream_conv2d_4_source_20_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_1 <= _source_stream_conv2d_4_source_20_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_2 <= _source_stream_conv2d_4_source_20_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_3 <= _source_stream_conv2d_4_source_20_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1031 <= _stream_conv2d_4_source_20_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_idle <= 0;
        _stream_conv2d_4_source_20_source_ram_raddr <= _stream_conv2d_4_source_20_source_pat_all_offset;
        _stream_conv2d_4_source_20_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= _source_stream_conv2d_4_source_20_pat_cur_offset_0 + _source_stream_conv2d_4_source_20_pat_stride_buf_0;
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= _source_stream_conv2d_4_source_20_pat_cur_offset_1 + _source_stream_conv2d_4_source_20_pat_stride_buf_1;
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= _source_stream_conv2d_4_source_20_pat_cur_offset_2 + _source_stream_conv2d_4_source_20_pat_stride_buf_2;
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= _source_stream_conv2d_4_source_20_pat_cur_offset_3 + _source_stream_conv2d_4_source_20_pat_stride_buf_3;
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_20_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_idle <= 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_idle <= 1;
      end 
      if(_set_flag_298) begin
        _stream_conv2d_4_source_21_source_mode <= 5'b10;
        _stream_conv2d_4_source_21_source_offset <= conv2d_4_stream_act_local_1 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_298) begin
        _source_stream_conv2d_4_source_21_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_298) begin
        _source_stream_conv2d_4_source_21_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_21_pat_stride_1 <= 0;
      end 
      if(_set_flag_298) begin
        _source_stream_conv2d_4_source_21_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_298) begin
        _source_stream_conv2d_4_source_21_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_298) begin
        _stream_conv2d_4_source_21_source_sel <= 4;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_offset_buf <= _stream_conv2d_4_source_21_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_0 <= _source_stream_conv2d_4_source_21_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_1 <= _source_stream_conv2d_4_source_21_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_2 <= _source_stream_conv2d_4_source_21_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_3 <= _source_stream_conv2d_4_source_21_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_0 <= _source_stream_conv2d_4_source_21_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_1 <= _source_stream_conv2d_4_source_21_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_2 <= _source_stream_conv2d_4_source_21_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_3 <= _source_stream_conv2d_4_source_21_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1032 <= _stream_conv2d_4_source_21_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_idle <= 0;
        _stream_conv2d_4_source_21_source_ram_raddr <= _stream_conv2d_4_source_21_source_pat_all_offset;
        _stream_conv2d_4_source_21_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= _source_stream_conv2d_4_source_21_pat_cur_offset_0 + _source_stream_conv2d_4_source_21_pat_stride_buf_0;
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= _source_stream_conv2d_4_source_21_pat_cur_offset_1 + _source_stream_conv2d_4_source_21_pat_stride_buf_1;
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= _source_stream_conv2d_4_source_21_pat_cur_offset_2 + _source_stream_conv2d_4_source_21_pat_stride_buf_2;
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= _source_stream_conv2d_4_source_21_pat_cur_offset_3 + _source_stream_conv2d_4_source_21_pat_stride_buf_3;
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_21_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_idle <= 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_idle <= 1;
      end 
      if(_set_flag_301) begin
        _stream_conv2d_4_source_22_source_mode <= 5'b10;
        _stream_conv2d_4_source_22_source_offset <= conv2d_4_stream_act_local_2 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_301) begin
        _source_stream_conv2d_4_source_22_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_301) begin
        _source_stream_conv2d_4_source_22_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_22_pat_stride_1 <= 0;
      end 
      if(_set_flag_301) begin
        _source_stream_conv2d_4_source_22_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_301) begin
        _source_stream_conv2d_4_source_22_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_301) begin
        _stream_conv2d_4_source_22_source_sel <= 5;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_offset_buf <= _stream_conv2d_4_source_22_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_0 <= _source_stream_conv2d_4_source_22_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_1 <= _source_stream_conv2d_4_source_22_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_2 <= _source_stream_conv2d_4_source_22_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_3 <= _source_stream_conv2d_4_source_22_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_0 <= _source_stream_conv2d_4_source_22_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_1 <= _source_stream_conv2d_4_source_22_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_2 <= _source_stream_conv2d_4_source_22_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_3 <= _source_stream_conv2d_4_source_22_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1033 <= _stream_conv2d_4_source_22_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_idle <= 0;
        _stream_conv2d_4_source_22_source_ram_raddr <= _stream_conv2d_4_source_22_source_pat_all_offset;
        _stream_conv2d_4_source_22_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= _source_stream_conv2d_4_source_22_pat_cur_offset_0 + _source_stream_conv2d_4_source_22_pat_stride_buf_0;
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= _source_stream_conv2d_4_source_22_pat_cur_offset_1 + _source_stream_conv2d_4_source_22_pat_stride_buf_1;
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= _source_stream_conv2d_4_source_22_pat_cur_offset_2 + _source_stream_conv2d_4_source_22_pat_stride_buf_2;
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= _source_stream_conv2d_4_source_22_pat_cur_offset_3 + _source_stream_conv2d_4_source_22_pat_stride_buf_3;
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_22_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_idle <= 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_idle <= 1;
      end 
      if(_set_flag_304) begin
        _stream_conv2d_4_source_23_source_mode <= 5'b10;
        _stream_conv2d_4_source_23_source_offset <= conv2d_4_stream_act_local_3 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_304) begin
        _source_stream_conv2d_4_source_23_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_23_pat_stride_0 <= 1;
      end 
      if(_set_flag_304) begin
        _source_stream_conv2d_4_source_23_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_23_pat_stride_1 <= 0;
      end 
      if(_set_flag_304) begin
        _source_stream_conv2d_4_source_23_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_23_pat_stride_2 <= 0;
      end 
      if(_set_flag_304) begin
        _source_stream_conv2d_4_source_23_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_23_pat_stride_3 <= 0;
      end 
      if(_set_flag_304) begin
        _stream_conv2d_4_source_23_source_sel <= 6;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_offset_buf <= _stream_conv2d_4_source_23_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_0 <= _source_stream_conv2d_4_source_23_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_1 <= _source_stream_conv2d_4_source_23_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_2 <= _source_stream_conv2d_4_source_23_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_3 <= _source_stream_conv2d_4_source_23_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_0 <= _source_stream_conv2d_4_source_23_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_1 <= _source_stream_conv2d_4_source_23_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_2 <= _source_stream_conv2d_4_source_23_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_3 <= _source_stream_conv2d_4_source_23_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1034 <= _stream_conv2d_4_source_23_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_idle <= 0;
        _stream_conv2d_4_source_23_source_ram_raddr <= _stream_conv2d_4_source_23_source_pat_all_offset;
        _stream_conv2d_4_source_23_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= _source_stream_conv2d_4_source_23_pat_cur_offset_0 + _source_stream_conv2d_4_source_23_pat_stride_buf_0;
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= _source_stream_conv2d_4_source_23_pat_cur_offset_1 + _source_stream_conv2d_4_source_23_pat_stride_buf_1;
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= _source_stream_conv2d_4_source_23_pat_cur_offset_2 + _source_stream_conv2d_4_source_23_pat_stride_buf_2;
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= _source_stream_conv2d_4_source_23_pat_cur_offset_3 + _source_stream_conv2d_4_source_23_pat_stride_buf_3;
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_23_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_idle <= 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_idle <= 1;
      end 
      if(_set_flag_307) begin
        _stream_conv2d_4_source_24_source_mode <= 5'b10;
        _stream_conv2d_4_source_24_source_offset <= conv2d_4_stream_act_local_4 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_307) begin
        _source_stream_conv2d_4_source_24_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_24_pat_stride_0 <= 1;
      end 
      if(_set_flag_307) begin
        _source_stream_conv2d_4_source_24_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_24_pat_stride_1 <= 0;
      end 
      if(_set_flag_307) begin
        _source_stream_conv2d_4_source_24_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_24_pat_stride_2 <= 0;
      end 
      if(_set_flag_307) begin
        _source_stream_conv2d_4_source_24_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_24_pat_stride_3 <= 0;
      end 
      if(_set_flag_307) begin
        _stream_conv2d_4_source_24_source_sel <= 7;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_offset_buf <= _stream_conv2d_4_source_24_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_0 <= _source_stream_conv2d_4_source_24_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_1 <= _source_stream_conv2d_4_source_24_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_2 <= _source_stream_conv2d_4_source_24_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_3 <= _source_stream_conv2d_4_source_24_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_0 <= _source_stream_conv2d_4_source_24_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_1 <= _source_stream_conv2d_4_source_24_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_2 <= _source_stream_conv2d_4_source_24_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_3 <= _source_stream_conv2d_4_source_24_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1035 <= _stream_conv2d_4_source_24_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_idle <= 0;
        _stream_conv2d_4_source_24_source_ram_raddr <= _stream_conv2d_4_source_24_source_pat_all_offset;
        _stream_conv2d_4_source_24_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= _source_stream_conv2d_4_source_24_pat_cur_offset_0 + _source_stream_conv2d_4_source_24_pat_stride_buf_0;
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= _source_stream_conv2d_4_source_24_pat_cur_offset_1 + _source_stream_conv2d_4_source_24_pat_stride_buf_1;
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= _source_stream_conv2d_4_source_24_pat_cur_offset_2 + _source_stream_conv2d_4_source_24_pat_stride_buf_2;
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= _source_stream_conv2d_4_source_24_pat_cur_offset_3 + _source_stream_conv2d_4_source_24_pat_stride_buf_3;
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_24_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_idle <= 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_idle <= 1;
      end 
      if(_set_flag_310) begin
        _stream_conv2d_4_source_25_source_mode <= 5'b10;
        _stream_conv2d_4_source_25_source_offset <= conv2d_4_stream_act_local_5 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_310) begin
        _source_stream_conv2d_4_source_25_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_25_pat_stride_0 <= 1;
      end 
      if(_set_flag_310) begin
        _source_stream_conv2d_4_source_25_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_25_pat_stride_1 <= 0;
      end 
      if(_set_flag_310) begin
        _source_stream_conv2d_4_source_25_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_25_pat_stride_2 <= 0;
      end 
      if(_set_flag_310) begin
        _source_stream_conv2d_4_source_25_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_25_pat_stride_3 <= 0;
      end 
      if(_set_flag_310) begin
        _stream_conv2d_4_source_25_source_sel <= 8;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_offset_buf <= _stream_conv2d_4_source_25_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_0 <= _source_stream_conv2d_4_source_25_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_1 <= _source_stream_conv2d_4_source_25_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_2 <= _source_stream_conv2d_4_source_25_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_3 <= _source_stream_conv2d_4_source_25_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_0 <= _source_stream_conv2d_4_source_25_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_1 <= _source_stream_conv2d_4_source_25_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_2 <= _source_stream_conv2d_4_source_25_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_3 <= _source_stream_conv2d_4_source_25_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1036 <= _stream_conv2d_4_source_25_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_idle <= 0;
        _stream_conv2d_4_source_25_source_ram_raddr <= _stream_conv2d_4_source_25_source_pat_all_offset;
        _stream_conv2d_4_source_25_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= _source_stream_conv2d_4_source_25_pat_cur_offset_0 + _source_stream_conv2d_4_source_25_pat_stride_buf_0;
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= _source_stream_conv2d_4_source_25_pat_cur_offset_1 + _source_stream_conv2d_4_source_25_pat_stride_buf_1;
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= _source_stream_conv2d_4_source_25_pat_cur_offset_2 + _source_stream_conv2d_4_source_25_pat_stride_buf_2;
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= _source_stream_conv2d_4_source_25_pat_cur_offset_3 + _source_stream_conv2d_4_source_25_pat_stride_buf_3;
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_25_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_idle <= 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_idle <= 1;
      end 
      if(_set_flag_313) begin
        _stream_conv2d_4_source_26_source_mode <= 5'b10;
        _stream_conv2d_4_source_26_source_offset <= conv2d_4_stream_act_local_6 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_313) begin
        _source_stream_conv2d_4_source_26_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_26_pat_stride_0 <= 1;
      end 
      if(_set_flag_313) begin
        _source_stream_conv2d_4_source_26_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_26_pat_stride_1 <= 0;
      end 
      if(_set_flag_313) begin
        _source_stream_conv2d_4_source_26_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_26_pat_stride_2 <= 0;
      end 
      if(_set_flag_313) begin
        _source_stream_conv2d_4_source_26_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_26_pat_stride_3 <= 0;
      end 
      if(_set_flag_313) begin
        _stream_conv2d_4_source_26_source_sel <= 9;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_offset_buf <= _stream_conv2d_4_source_26_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_0 <= _source_stream_conv2d_4_source_26_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_1 <= _source_stream_conv2d_4_source_26_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_2 <= _source_stream_conv2d_4_source_26_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_3 <= _source_stream_conv2d_4_source_26_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_0 <= _source_stream_conv2d_4_source_26_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_1 <= _source_stream_conv2d_4_source_26_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_2 <= _source_stream_conv2d_4_source_26_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_3 <= _source_stream_conv2d_4_source_26_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1037 <= _stream_conv2d_4_source_26_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_idle <= 0;
        _stream_conv2d_4_source_26_source_ram_raddr <= _stream_conv2d_4_source_26_source_pat_all_offset;
        _stream_conv2d_4_source_26_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= _source_stream_conv2d_4_source_26_pat_cur_offset_0 + _source_stream_conv2d_4_source_26_pat_stride_buf_0;
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= _source_stream_conv2d_4_source_26_pat_cur_offset_1 + _source_stream_conv2d_4_source_26_pat_stride_buf_1;
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= _source_stream_conv2d_4_source_26_pat_cur_offset_2 + _source_stream_conv2d_4_source_26_pat_stride_buf_2;
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= _source_stream_conv2d_4_source_26_pat_cur_offset_3 + _source_stream_conv2d_4_source_26_pat_stride_buf_3;
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_26_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_idle <= 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_idle <= 1;
      end 
      if(_set_flag_316) begin
        _stream_conv2d_4_source_27_source_mode <= 5'b10;
        _stream_conv2d_4_source_27_source_offset <= conv2d_4_stream_act_local_7 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_316) begin
        _source_stream_conv2d_4_source_27_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_27_pat_stride_0 <= 1;
      end 
      if(_set_flag_316) begin
        _source_stream_conv2d_4_source_27_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_27_pat_stride_1 <= 0;
      end 
      if(_set_flag_316) begin
        _source_stream_conv2d_4_source_27_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_27_pat_stride_2 <= 0;
      end 
      if(_set_flag_316) begin
        _source_stream_conv2d_4_source_27_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_27_pat_stride_3 <= 0;
      end 
      if(_set_flag_316) begin
        _stream_conv2d_4_source_27_source_sel <= 10;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_offset_buf <= _stream_conv2d_4_source_27_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_0 <= _source_stream_conv2d_4_source_27_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_1 <= _source_stream_conv2d_4_source_27_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_2 <= _source_stream_conv2d_4_source_27_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_3 <= _source_stream_conv2d_4_source_27_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_0 <= _source_stream_conv2d_4_source_27_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_1 <= _source_stream_conv2d_4_source_27_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_2 <= _source_stream_conv2d_4_source_27_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_3 <= _source_stream_conv2d_4_source_27_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1038 <= _stream_conv2d_4_source_27_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_idle <= 0;
        _stream_conv2d_4_source_27_source_ram_raddr <= _stream_conv2d_4_source_27_source_pat_all_offset;
        _stream_conv2d_4_source_27_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= _source_stream_conv2d_4_source_27_pat_cur_offset_0 + _source_stream_conv2d_4_source_27_pat_stride_buf_0;
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= _source_stream_conv2d_4_source_27_pat_cur_offset_1 + _source_stream_conv2d_4_source_27_pat_stride_buf_1;
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= _source_stream_conv2d_4_source_27_pat_cur_offset_2 + _source_stream_conv2d_4_source_27_pat_stride_buf_2;
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= _source_stream_conv2d_4_source_27_pat_cur_offset_3 + _source_stream_conv2d_4_source_27_pat_stride_buf_3;
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_27_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_idle <= 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_idle <= 1;
      end 
      if(_set_flag_319) begin
        _stream_conv2d_4_source_28_source_mode <= 5'b10;
        _stream_conv2d_4_source_28_source_offset <= conv2d_4_stream_act_local_8 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_319) begin
        _source_stream_conv2d_4_source_28_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_28_pat_stride_0 <= 1;
      end 
      if(_set_flag_319) begin
        _source_stream_conv2d_4_source_28_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_28_pat_stride_1 <= 0;
      end 
      if(_set_flag_319) begin
        _source_stream_conv2d_4_source_28_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_28_pat_stride_2 <= 0;
      end 
      if(_set_flag_319) begin
        _source_stream_conv2d_4_source_28_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_28_pat_stride_3 <= 0;
      end 
      if(_set_flag_319) begin
        _stream_conv2d_4_source_28_source_sel <= 11;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_offset_buf <= _stream_conv2d_4_source_28_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_0 <= _source_stream_conv2d_4_source_28_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_1 <= _source_stream_conv2d_4_source_28_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_2 <= _source_stream_conv2d_4_source_28_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_3 <= _source_stream_conv2d_4_source_28_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_0 <= _source_stream_conv2d_4_source_28_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_1 <= _source_stream_conv2d_4_source_28_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_2 <= _source_stream_conv2d_4_source_28_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_3 <= _source_stream_conv2d_4_source_28_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1039 <= _stream_conv2d_4_source_28_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_idle <= 0;
        _stream_conv2d_4_source_28_source_ram_raddr <= _stream_conv2d_4_source_28_source_pat_all_offset;
        _stream_conv2d_4_source_28_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= _source_stream_conv2d_4_source_28_pat_cur_offset_0 + _source_stream_conv2d_4_source_28_pat_stride_buf_0;
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= _source_stream_conv2d_4_source_28_pat_cur_offset_1 + _source_stream_conv2d_4_source_28_pat_stride_buf_1;
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= _source_stream_conv2d_4_source_28_pat_cur_offset_2 + _source_stream_conv2d_4_source_28_pat_stride_buf_2;
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= _source_stream_conv2d_4_source_28_pat_cur_offset_3 + _source_stream_conv2d_4_source_28_pat_stride_buf_3;
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_28_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_idle <= 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_idle <= 1;
      end 
      if(_set_flag_322) begin
        _stream_conv2d_4_source_29_source_mode <= 5'b10;
        _stream_conv2d_4_source_29_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_322) begin
        _source_stream_conv2d_4_source_29_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_29_pat_stride_0 <= 1;
      end 
      if(_set_flag_322) begin
        _source_stream_conv2d_4_source_29_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_29_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_322) begin
        _source_stream_conv2d_4_source_29_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_29_pat_stride_2 <= 0;
      end 
      if(_set_flag_322) begin
        _source_stream_conv2d_4_source_29_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_29_pat_stride_3 <= 0;
      end 
      if(_set_flag_322) begin
        _stream_conv2d_4_source_29_source_sel <= 12;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_offset_buf <= _stream_conv2d_4_source_29_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_0 <= _source_stream_conv2d_4_source_29_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_1 <= _source_stream_conv2d_4_source_29_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_2 <= _source_stream_conv2d_4_source_29_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_3 <= _source_stream_conv2d_4_source_29_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_0 <= _source_stream_conv2d_4_source_29_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_1 <= _source_stream_conv2d_4_source_29_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_2 <= _source_stream_conv2d_4_source_29_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_3 <= _source_stream_conv2d_4_source_29_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1328 <= _stream_conv2d_4_source_29_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_idle <= 0;
        _stream_conv2d_4_source_29_source_ram_raddr <= _stream_conv2d_4_source_29_source_pat_all_offset;
        _stream_conv2d_4_source_29_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= _source_stream_conv2d_4_source_29_pat_cur_offset_0 + _source_stream_conv2d_4_source_29_pat_stride_buf_0;
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= _source_stream_conv2d_4_source_29_pat_cur_offset_1 + _source_stream_conv2d_4_source_29_pat_stride_buf_1;
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= _source_stream_conv2d_4_source_29_pat_cur_offset_2 + _source_stream_conv2d_4_source_29_pat_stride_buf_2;
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= _source_stream_conv2d_4_source_29_pat_cur_offset_3 + _source_stream_conv2d_4_source_29_pat_stride_buf_3;
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_29_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_idle <= 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_idle <= 1;
      end 
      if(_set_flag_325) begin
        _stream_conv2d_4_source_30_source_mode <= 5'b10;
        _stream_conv2d_4_source_30_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_325) begin
        _source_stream_conv2d_4_source_30_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_30_pat_stride_0 <= 1;
      end 
      if(_set_flag_325) begin
        _source_stream_conv2d_4_source_30_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_30_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_325) begin
        _source_stream_conv2d_4_source_30_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_30_pat_stride_2 <= 0;
      end 
      if(_set_flag_325) begin
        _source_stream_conv2d_4_source_30_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_30_pat_stride_3 <= 0;
      end 
      if(_set_flag_325) begin
        _stream_conv2d_4_source_30_source_sel <= 13;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_offset_buf <= _stream_conv2d_4_source_30_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_0 <= _source_stream_conv2d_4_source_30_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_1 <= _source_stream_conv2d_4_source_30_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_2 <= _source_stream_conv2d_4_source_30_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_3 <= _source_stream_conv2d_4_source_30_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_0 <= _source_stream_conv2d_4_source_30_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_1 <= _source_stream_conv2d_4_source_30_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_2 <= _source_stream_conv2d_4_source_30_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_3 <= _source_stream_conv2d_4_source_30_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1329 <= _stream_conv2d_4_source_30_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_idle <= 0;
        _stream_conv2d_4_source_30_source_ram_raddr <= _stream_conv2d_4_source_30_source_pat_all_offset;
        _stream_conv2d_4_source_30_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= _source_stream_conv2d_4_source_30_pat_cur_offset_0 + _source_stream_conv2d_4_source_30_pat_stride_buf_0;
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= _source_stream_conv2d_4_source_30_pat_cur_offset_1 + _source_stream_conv2d_4_source_30_pat_stride_buf_1;
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= _source_stream_conv2d_4_source_30_pat_cur_offset_2 + _source_stream_conv2d_4_source_30_pat_stride_buf_2;
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= _source_stream_conv2d_4_source_30_pat_cur_offset_3 + _source_stream_conv2d_4_source_30_pat_stride_buf_3;
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_30_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_idle <= 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_idle <= 1;
      end 
      if(_set_flag_328) begin
        _stream_conv2d_4_source_31_source_mode <= 5'b10;
        _stream_conv2d_4_source_31_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_328) begin
        _source_stream_conv2d_4_source_31_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_31_pat_stride_0 <= 1;
      end 
      if(_set_flag_328) begin
        _source_stream_conv2d_4_source_31_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_31_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_328) begin
        _source_stream_conv2d_4_source_31_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_31_pat_stride_2 <= 0;
      end 
      if(_set_flag_328) begin
        _source_stream_conv2d_4_source_31_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_31_pat_stride_3 <= 0;
      end 
      if(_set_flag_328) begin
        _stream_conv2d_4_source_31_source_sel <= 14;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_offset_buf <= _stream_conv2d_4_source_31_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_0 <= _source_stream_conv2d_4_source_31_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_1 <= _source_stream_conv2d_4_source_31_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_2 <= _source_stream_conv2d_4_source_31_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_3 <= _source_stream_conv2d_4_source_31_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_0 <= _source_stream_conv2d_4_source_31_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_1 <= _source_stream_conv2d_4_source_31_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_2 <= _source_stream_conv2d_4_source_31_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_3 <= _source_stream_conv2d_4_source_31_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1330 <= _stream_conv2d_4_source_31_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_idle <= 0;
        _stream_conv2d_4_source_31_source_ram_raddr <= _stream_conv2d_4_source_31_source_pat_all_offset;
        _stream_conv2d_4_source_31_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= _source_stream_conv2d_4_source_31_pat_cur_offset_0 + _source_stream_conv2d_4_source_31_pat_stride_buf_0;
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= _source_stream_conv2d_4_source_31_pat_cur_offset_1 + _source_stream_conv2d_4_source_31_pat_stride_buf_1;
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= _source_stream_conv2d_4_source_31_pat_cur_offset_2 + _source_stream_conv2d_4_source_31_pat_stride_buf_2;
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= _source_stream_conv2d_4_source_31_pat_cur_offset_3 + _source_stream_conv2d_4_source_31_pat_stride_buf_3;
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_31_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_idle <= 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_idle <= 1;
      end 
      if(_set_flag_331) begin
        _stream_conv2d_4_source_32_source_mode <= 5'b10;
        _stream_conv2d_4_source_32_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_331) begin
        _source_stream_conv2d_4_source_32_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_32_pat_stride_0 <= 1;
      end 
      if(_set_flag_331) begin
        _source_stream_conv2d_4_source_32_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_32_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_331) begin
        _source_stream_conv2d_4_source_32_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_32_pat_stride_2 <= 0;
      end 
      if(_set_flag_331) begin
        _source_stream_conv2d_4_source_32_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_32_pat_stride_3 <= 0;
      end 
      if(_set_flag_331) begin
        _stream_conv2d_4_source_32_source_sel <= 15;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_offset_buf <= _stream_conv2d_4_source_32_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_0 <= _source_stream_conv2d_4_source_32_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_1 <= _source_stream_conv2d_4_source_32_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_2 <= _source_stream_conv2d_4_source_32_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_3 <= _source_stream_conv2d_4_source_32_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_0 <= _source_stream_conv2d_4_source_32_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_1 <= _source_stream_conv2d_4_source_32_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_2 <= _source_stream_conv2d_4_source_32_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_3 <= _source_stream_conv2d_4_source_32_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1331 <= _stream_conv2d_4_source_32_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_idle <= 0;
        _stream_conv2d_4_source_32_source_ram_raddr <= _stream_conv2d_4_source_32_source_pat_all_offset;
        _stream_conv2d_4_source_32_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= _source_stream_conv2d_4_source_32_pat_cur_offset_0 + _source_stream_conv2d_4_source_32_pat_stride_buf_0;
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= _source_stream_conv2d_4_source_32_pat_cur_offset_1 + _source_stream_conv2d_4_source_32_pat_stride_buf_1;
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= _source_stream_conv2d_4_source_32_pat_cur_offset_2 + _source_stream_conv2d_4_source_32_pat_stride_buf_2;
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= _source_stream_conv2d_4_source_32_pat_cur_offset_3 + _source_stream_conv2d_4_source_32_pat_stride_buf_3;
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_32_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_idle <= 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_idle <= 1;
      end 
      if(_set_flag_334) begin
        _stream_conv2d_4_source_33_source_mode <= 5'b10;
        _stream_conv2d_4_source_33_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_33_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_33_pat_stride_0 <= 1;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_33_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_33_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_33_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_33_pat_stride_2 <= 0;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_33_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_33_pat_stride_3 <= 0;
      end 
      if(_set_flag_334) begin
        _stream_conv2d_4_source_33_source_sel <= 16;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_offset_buf <= _stream_conv2d_4_source_33_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_0 <= _source_stream_conv2d_4_source_33_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_1 <= _source_stream_conv2d_4_source_33_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_2 <= _source_stream_conv2d_4_source_33_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_3 <= _source_stream_conv2d_4_source_33_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_0 <= _source_stream_conv2d_4_source_33_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_1 <= _source_stream_conv2d_4_source_33_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_2 <= _source_stream_conv2d_4_source_33_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_3 <= _source_stream_conv2d_4_source_33_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1332 <= _stream_conv2d_4_source_33_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_idle <= 0;
        _stream_conv2d_4_source_33_source_ram_raddr <= _stream_conv2d_4_source_33_source_pat_all_offset;
        _stream_conv2d_4_source_33_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= _source_stream_conv2d_4_source_33_pat_cur_offset_0 + _source_stream_conv2d_4_source_33_pat_stride_buf_0;
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= _source_stream_conv2d_4_source_33_pat_cur_offset_1 + _source_stream_conv2d_4_source_33_pat_stride_buf_1;
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= _source_stream_conv2d_4_source_33_pat_cur_offset_2 + _source_stream_conv2d_4_source_33_pat_stride_buf_2;
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= _source_stream_conv2d_4_source_33_pat_cur_offset_3 + _source_stream_conv2d_4_source_33_pat_stride_buf_3;
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_33_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_idle <= 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_idle <= 1;
      end 
      if(_set_flag_337) begin
        _stream_conv2d_4_source_34_source_mode <= 5'b10;
        _stream_conv2d_4_source_34_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_337) begin
        _source_stream_conv2d_4_source_34_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_34_pat_stride_0 <= 1;
      end 
      if(_set_flag_337) begin
        _source_stream_conv2d_4_source_34_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_34_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_337) begin
        _source_stream_conv2d_4_source_34_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_34_pat_stride_2 <= 0;
      end 
      if(_set_flag_337) begin
        _source_stream_conv2d_4_source_34_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_34_pat_stride_3 <= 0;
      end 
      if(_set_flag_337) begin
        _stream_conv2d_4_source_34_source_sel <= 17;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_offset_buf <= _stream_conv2d_4_source_34_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_0 <= _source_stream_conv2d_4_source_34_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_1 <= _source_stream_conv2d_4_source_34_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_2 <= _source_stream_conv2d_4_source_34_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_3 <= _source_stream_conv2d_4_source_34_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_0 <= _source_stream_conv2d_4_source_34_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_1 <= _source_stream_conv2d_4_source_34_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_2 <= _source_stream_conv2d_4_source_34_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_3 <= _source_stream_conv2d_4_source_34_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1333 <= _stream_conv2d_4_source_34_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_idle <= 0;
        _stream_conv2d_4_source_34_source_ram_raddr <= _stream_conv2d_4_source_34_source_pat_all_offset;
        _stream_conv2d_4_source_34_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= _source_stream_conv2d_4_source_34_pat_cur_offset_0 + _source_stream_conv2d_4_source_34_pat_stride_buf_0;
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= _source_stream_conv2d_4_source_34_pat_cur_offset_1 + _source_stream_conv2d_4_source_34_pat_stride_buf_1;
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= _source_stream_conv2d_4_source_34_pat_cur_offset_2 + _source_stream_conv2d_4_source_34_pat_stride_buf_2;
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= _source_stream_conv2d_4_source_34_pat_cur_offset_3 + _source_stream_conv2d_4_source_34_pat_stride_buf_3;
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_34_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_idle <= 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_idle <= 1;
      end 
      if(_set_flag_340) begin
        _stream_conv2d_4_source_35_source_mode <= 5'b10;
        _stream_conv2d_4_source_35_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_340) begin
        _source_stream_conv2d_4_source_35_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_35_pat_stride_0 <= 1;
      end 
      if(_set_flag_340) begin
        _source_stream_conv2d_4_source_35_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_35_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_340) begin
        _source_stream_conv2d_4_source_35_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_35_pat_stride_2 <= 0;
      end 
      if(_set_flag_340) begin
        _source_stream_conv2d_4_source_35_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_35_pat_stride_3 <= 0;
      end 
      if(_set_flag_340) begin
        _stream_conv2d_4_source_35_source_sel <= 18;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_offset_buf <= _stream_conv2d_4_source_35_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_0 <= _source_stream_conv2d_4_source_35_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_1 <= _source_stream_conv2d_4_source_35_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_2 <= _source_stream_conv2d_4_source_35_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_3 <= _source_stream_conv2d_4_source_35_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_0 <= _source_stream_conv2d_4_source_35_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_1 <= _source_stream_conv2d_4_source_35_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_2 <= _source_stream_conv2d_4_source_35_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_3 <= _source_stream_conv2d_4_source_35_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1334 <= _stream_conv2d_4_source_35_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_idle <= 0;
        _stream_conv2d_4_source_35_source_ram_raddr <= _stream_conv2d_4_source_35_source_pat_all_offset;
        _stream_conv2d_4_source_35_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= _source_stream_conv2d_4_source_35_pat_cur_offset_0 + _source_stream_conv2d_4_source_35_pat_stride_buf_0;
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= _source_stream_conv2d_4_source_35_pat_cur_offset_1 + _source_stream_conv2d_4_source_35_pat_stride_buf_1;
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= _source_stream_conv2d_4_source_35_pat_cur_offset_2 + _source_stream_conv2d_4_source_35_pat_stride_buf_2;
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= _source_stream_conv2d_4_source_35_pat_cur_offset_3 + _source_stream_conv2d_4_source_35_pat_stride_buf_3;
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_35_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_idle <= 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_idle <= 1;
      end 
      if(_set_flag_343) begin
        _stream_conv2d_4_source_36_source_mode <= 5'b10;
        _stream_conv2d_4_source_36_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_343) begin
        _source_stream_conv2d_4_source_36_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_36_pat_stride_0 <= 1;
      end 
      if(_set_flag_343) begin
        _source_stream_conv2d_4_source_36_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_36_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_343) begin
        _source_stream_conv2d_4_source_36_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_36_pat_stride_2 <= 0;
      end 
      if(_set_flag_343) begin
        _source_stream_conv2d_4_source_36_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_36_pat_stride_3 <= 0;
      end 
      if(_set_flag_343) begin
        _stream_conv2d_4_source_36_source_sel <= 19;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_offset_buf <= _stream_conv2d_4_source_36_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_0 <= _source_stream_conv2d_4_source_36_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_1 <= _source_stream_conv2d_4_source_36_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_2 <= _source_stream_conv2d_4_source_36_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_3 <= _source_stream_conv2d_4_source_36_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_0 <= _source_stream_conv2d_4_source_36_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_1 <= _source_stream_conv2d_4_source_36_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_2 <= _source_stream_conv2d_4_source_36_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_3 <= _source_stream_conv2d_4_source_36_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1335 <= _stream_conv2d_4_source_36_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_idle <= 0;
        _stream_conv2d_4_source_36_source_ram_raddr <= _stream_conv2d_4_source_36_source_pat_all_offset;
        _stream_conv2d_4_source_36_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= _source_stream_conv2d_4_source_36_pat_cur_offset_0 + _source_stream_conv2d_4_source_36_pat_stride_buf_0;
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= _source_stream_conv2d_4_source_36_pat_cur_offset_1 + _source_stream_conv2d_4_source_36_pat_stride_buf_1;
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= _source_stream_conv2d_4_source_36_pat_cur_offset_2 + _source_stream_conv2d_4_source_36_pat_stride_buf_2;
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= _source_stream_conv2d_4_source_36_pat_cur_offset_3 + _source_stream_conv2d_4_source_36_pat_stride_buf_3;
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_36_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_idle <= 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_idle <= 1;
      end 
      if(_set_flag_346) begin
        _stream_conv2d_4_source_37_source_mode <= 5'b10;
        _stream_conv2d_4_source_37_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_346) begin
        _source_stream_conv2d_4_source_37_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_37_pat_stride_0 <= 1;
      end 
      if(_set_flag_346) begin
        _source_stream_conv2d_4_source_37_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_37_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_346) begin
        _source_stream_conv2d_4_source_37_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_37_pat_stride_2 <= 0;
      end 
      if(_set_flag_346) begin
        _source_stream_conv2d_4_source_37_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_37_pat_stride_3 <= 0;
      end 
      if(_set_flag_346) begin
        _stream_conv2d_4_source_37_source_sel <= 20;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_offset_buf <= _stream_conv2d_4_source_37_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_0 <= _source_stream_conv2d_4_source_37_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_1 <= _source_stream_conv2d_4_source_37_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_2 <= _source_stream_conv2d_4_source_37_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_3 <= _source_stream_conv2d_4_source_37_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_0 <= _source_stream_conv2d_4_source_37_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_1 <= _source_stream_conv2d_4_source_37_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_2 <= _source_stream_conv2d_4_source_37_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_3 <= _source_stream_conv2d_4_source_37_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1336 <= _stream_conv2d_4_source_37_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_idle <= 0;
        _stream_conv2d_4_source_37_source_ram_raddr <= _stream_conv2d_4_source_37_source_pat_all_offset;
        _stream_conv2d_4_source_37_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= _source_stream_conv2d_4_source_37_pat_cur_offset_0 + _source_stream_conv2d_4_source_37_pat_stride_buf_0;
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= _source_stream_conv2d_4_source_37_pat_cur_offset_1 + _source_stream_conv2d_4_source_37_pat_stride_buf_1;
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= _source_stream_conv2d_4_source_37_pat_cur_offset_2 + _source_stream_conv2d_4_source_37_pat_stride_buf_2;
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= _source_stream_conv2d_4_source_37_pat_cur_offset_3 + _source_stream_conv2d_4_source_37_pat_stride_buf_3;
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_37_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_idle <= 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_idle <= 1;
      end 
      if(_set_flag_349) begin
        _stream_conv2d_4_source_38_source_mode <= 5'b10;
        _stream_conv2d_4_source_38_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_349) begin
        _source_stream_conv2d_4_source_38_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_38_pat_stride_0 <= 1;
      end 
      if(_set_flag_349) begin
        _source_stream_conv2d_4_source_38_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_38_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_349) begin
        _source_stream_conv2d_4_source_38_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_38_pat_stride_2 <= 0;
      end 
      if(_set_flag_349) begin
        _source_stream_conv2d_4_source_38_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_38_pat_stride_3 <= 0;
      end 
      if(_set_flag_349) begin
        _stream_conv2d_4_source_38_source_sel <= 21;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_38_source_offset_buf <= _stream_conv2d_4_source_38_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_count_0 <= _source_stream_conv2d_4_source_38_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_count_1 <= _source_stream_conv2d_4_source_38_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_count_2 <= _source_stream_conv2d_4_source_38_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_count_3 <= _source_stream_conv2d_4_source_38_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_size_buf_0 <= _source_stream_conv2d_4_source_38_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_size_buf_1 <= _source_stream_conv2d_4_source_38_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_size_buf_2 <= _source_stream_conv2d_4_source_38_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_size_buf_3 <= _source_stream_conv2d_4_source_38_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_stride_buf_0 <= _source_stream_conv2d_4_source_38_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_stride_buf_1 <= _source_stream_conv2d_4_source_38_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_stride_buf_2 <= _source_stream_conv2d_4_source_38_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_stride_buf_3 <= _source_stream_conv2d_4_source_38_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1337 <= _stream_conv2d_4_source_38_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_38_idle <= 0;
        _stream_conv2d_4_source_38_source_ram_raddr <= _stream_conv2d_4_source_38_source_pat_all_offset;
        _stream_conv2d_4_source_38_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_0 <= _source_stream_conv2d_4_source_38_pat_cur_offset_0 + _source_stream_conv2d_4_source_38_pat_stride_buf_0;
        _source_stream_conv2d_4_source_38_pat_count_0 <= _source_stream_conv2d_4_source_38_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && (_source_stream_conv2d_4_source_38_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_38_pat_count_0 <= _source_stream_conv2d_4_source_38_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && (_source_stream_conv2d_4_source_38_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_1 <= _source_stream_conv2d_4_source_38_pat_cur_offset_1 + _source_stream_conv2d_4_source_38_pat_stride_buf_1;
        _source_stream_conv2d_4_source_38_pat_count_1 <= _source_stream_conv2d_4_source_38_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && (_source_stream_conv2d_4_source_38_pat_count_0 == 0) && (_source_stream_conv2d_4_source_38_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_38_pat_count_1 <= _source_stream_conv2d_4_source_38_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && ((_source_stream_conv2d_4_source_38_pat_count_0 == 0) && (_source_stream_conv2d_4_source_38_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_2 <= _source_stream_conv2d_4_source_38_pat_cur_offset_2 + _source_stream_conv2d_4_source_38_pat_stride_buf_2;
        _source_stream_conv2d_4_source_38_pat_count_2 <= _source_stream_conv2d_4_source_38_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && ((_source_stream_conv2d_4_source_38_pat_count_0 == 0) && (_source_stream_conv2d_4_source_38_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_38_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_38_pat_count_2 <= _source_stream_conv2d_4_source_38_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && ((_source_stream_conv2d_4_source_38_pat_count_0 == 0) && (_source_stream_conv2d_4_source_38_pat_count_1 == 0) && (_source_stream_conv2d_4_source_38_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_3 <= _source_stream_conv2d_4_source_38_pat_cur_offset_3 + _source_stream_conv2d_4_source_38_pat_stride_buf_3;
        _source_stream_conv2d_4_source_38_pat_count_3 <= _source_stream_conv2d_4_source_38_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && ((_source_stream_conv2d_4_source_38_pat_count_0 == 0) && (_source_stream_conv2d_4_source_38_pat_count_1 == 0) && (_source_stream_conv2d_4_source_38_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_38_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_38_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_38_pat_count_3 <= _source_stream_conv2d_4_source_38_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_38_source_ram_renable <= 0;
        _stream_conv2d_4_source_38_idle <= 1;
      end 
      if((_stream_conv2d_4_source_38_source_pat_fsm_20 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_38_source_ram_renable <= 0;
        _stream_conv2d_4_source_38_idle <= 1;
      end 
      if(_set_flag_352) begin
        _stream_conv2d_4_source_39_source_mode <= 5'b10;
        _stream_conv2d_4_source_39_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_352) begin
        _source_stream_conv2d_4_source_39_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_39_pat_stride_0 <= 1;
      end 
      if(_set_flag_352) begin
        _source_stream_conv2d_4_source_39_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_39_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_352) begin
        _source_stream_conv2d_4_source_39_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_39_pat_stride_2 <= 0;
      end 
      if(_set_flag_352) begin
        _source_stream_conv2d_4_source_39_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_39_pat_stride_3 <= 0;
      end 
      if(_set_flag_352) begin
        _stream_conv2d_4_source_39_source_sel <= 22;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_39_source_offset_buf <= _stream_conv2d_4_source_39_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_count_0 <= _source_stream_conv2d_4_source_39_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_count_1 <= _source_stream_conv2d_4_source_39_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_count_2 <= _source_stream_conv2d_4_source_39_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_count_3 <= _source_stream_conv2d_4_source_39_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_size_buf_0 <= _source_stream_conv2d_4_source_39_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_size_buf_1 <= _source_stream_conv2d_4_source_39_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_size_buf_2 <= _source_stream_conv2d_4_source_39_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_size_buf_3 <= _source_stream_conv2d_4_source_39_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_stride_buf_0 <= _source_stream_conv2d_4_source_39_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_stride_buf_1 <= _source_stream_conv2d_4_source_39_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_stride_buf_2 <= _source_stream_conv2d_4_source_39_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_stride_buf_3 <= _source_stream_conv2d_4_source_39_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1338 <= _stream_conv2d_4_source_39_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_39_idle <= 0;
        _stream_conv2d_4_source_39_source_ram_raddr <= _stream_conv2d_4_source_39_source_pat_all_offset;
        _stream_conv2d_4_source_39_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_0 <= _source_stream_conv2d_4_source_39_pat_cur_offset_0 + _source_stream_conv2d_4_source_39_pat_stride_buf_0;
        _source_stream_conv2d_4_source_39_pat_count_0 <= _source_stream_conv2d_4_source_39_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && (_source_stream_conv2d_4_source_39_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_39_pat_count_0 <= _source_stream_conv2d_4_source_39_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && (_source_stream_conv2d_4_source_39_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_1 <= _source_stream_conv2d_4_source_39_pat_cur_offset_1 + _source_stream_conv2d_4_source_39_pat_stride_buf_1;
        _source_stream_conv2d_4_source_39_pat_count_1 <= _source_stream_conv2d_4_source_39_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && (_source_stream_conv2d_4_source_39_pat_count_0 == 0) && (_source_stream_conv2d_4_source_39_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_39_pat_count_1 <= _source_stream_conv2d_4_source_39_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && ((_source_stream_conv2d_4_source_39_pat_count_0 == 0) && (_source_stream_conv2d_4_source_39_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_2 <= _source_stream_conv2d_4_source_39_pat_cur_offset_2 + _source_stream_conv2d_4_source_39_pat_stride_buf_2;
        _source_stream_conv2d_4_source_39_pat_count_2 <= _source_stream_conv2d_4_source_39_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && ((_source_stream_conv2d_4_source_39_pat_count_0 == 0) && (_source_stream_conv2d_4_source_39_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_39_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_39_pat_count_2 <= _source_stream_conv2d_4_source_39_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && ((_source_stream_conv2d_4_source_39_pat_count_0 == 0) && (_source_stream_conv2d_4_source_39_pat_count_1 == 0) && (_source_stream_conv2d_4_source_39_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_3 <= _source_stream_conv2d_4_source_39_pat_cur_offset_3 + _source_stream_conv2d_4_source_39_pat_stride_buf_3;
        _source_stream_conv2d_4_source_39_pat_count_3 <= _source_stream_conv2d_4_source_39_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && ((_source_stream_conv2d_4_source_39_pat_count_0 == 0) && (_source_stream_conv2d_4_source_39_pat_count_1 == 0) && (_source_stream_conv2d_4_source_39_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_39_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_39_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_39_pat_count_3 <= _source_stream_conv2d_4_source_39_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_39_source_ram_renable <= 0;
        _stream_conv2d_4_source_39_idle <= 1;
      end 
      if((_stream_conv2d_4_source_39_source_pat_fsm_21 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_39_source_ram_renable <= 0;
        _stream_conv2d_4_source_39_idle <= 1;
      end 
      if(_set_flag_355) begin
        _stream_conv2d_4_source_40_source_mode <= 5'b10;
        _stream_conv2d_4_source_40_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_355) begin
        _source_stream_conv2d_4_source_40_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_40_pat_stride_0 <= 1;
      end 
      if(_set_flag_355) begin
        _source_stream_conv2d_4_source_40_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_40_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_355) begin
        _source_stream_conv2d_4_source_40_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_40_pat_stride_2 <= 0;
      end 
      if(_set_flag_355) begin
        _source_stream_conv2d_4_source_40_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_40_pat_stride_3 <= 0;
      end 
      if(_set_flag_355) begin
        _stream_conv2d_4_source_40_source_sel <= 23;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_40_source_offset_buf <= _stream_conv2d_4_source_40_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_count_0 <= _source_stream_conv2d_4_source_40_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_count_1 <= _source_stream_conv2d_4_source_40_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_count_2 <= _source_stream_conv2d_4_source_40_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_count_3 <= _source_stream_conv2d_4_source_40_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_size_buf_0 <= _source_stream_conv2d_4_source_40_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_size_buf_1 <= _source_stream_conv2d_4_source_40_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_size_buf_2 <= _source_stream_conv2d_4_source_40_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_size_buf_3 <= _source_stream_conv2d_4_source_40_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_stride_buf_0 <= _source_stream_conv2d_4_source_40_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_stride_buf_1 <= _source_stream_conv2d_4_source_40_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_stride_buf_2 <= _source_stream_conv2d_4_source_40_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_stride_buf_3 <= _source_stream_conv2d_4_source_40_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1339 <= _stream_conv2d_4_source_40_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_40_idle <= 0;
        _stream_conv2d_4_source_40_source_ram_raddr <= _stream_conv2d_4_source_40_source_pat_all_offset;
        _stream_conv2d_4_source_40_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_0 <= _source_stream_conv2d_4_source_40_pat_cur_offset_0 + _source_stream_conv2d_4_source_40_pat_stride_buf_0;
        _source_stream_conv2d_4_source_40_pat_count_0 <= _source_stream_conv2d_4_source_40_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && (_source_stream_conv2d_4_source_40_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_40_pat_count_0 <= _source_stream_conv2d_4_source_40_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && (_source_stream_conv2d_4_source_40_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_1 <= _source_stream_conv2d_4_source_40_pat_cur_offset_1 + _source_stream_conv2d_4_source_40_pat_stride_buf_1;
        _source_stream_conv2d_4_source_40_pat_count_1 <= _source_stream_conv2d_4_source_40_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && (_source_stream_conv2d_4_source_40_pat_count_0 == 0) && (_source_stream_conv2d_4_source_40_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_40_pat_count_1 <= _source_stream_conv2d_4_source_40_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && ((_source_stream_conv2d_4_source_40_pat_count_0 == 0) && (_source_stream_conv2d_4_source_40_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_2 <= _source_stream_conv2d_4_source_40_pat_cur_offset_2 + _source_stream_conv2d_4_source_40_pat_stride_buf_2;
        _source_stream_conv2d_4_source_40_pat_count_2 <= _source_stream_conv2d_4_source_40_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && ((_source_stream_conv2d_4_source_40_pat_count_0 == 0) && (_source_stream_conv2d_4_source_40_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_40_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_40_pat_count_2 <= _source_stream_conv2d_4_source_40_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && ((_source_stream_conv2d_4_source_40_pat_count_0 == 0) && (_source_stream_conv2d_4_source_40_pat_count_1 == 0) && (_source_stream_conv2d_4_source_40_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_3 <= _source_stream_conv2d_4_source_40_pat_cur_offset_3 + _source_stream_conv2d_4_source_40_pat_stride_buf_3;
        _source_stream_conv2d_4_source_40_pat_count_3 <= _source_stream_conv2d_4_source_40_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && ((_source_stream_conv2d_4_source_40_pat_count_0 == 0) && (_source_stream_conv2d_4_source_40_pat_count_1 == 0) && (_source_stream_conv2d_4_source_40_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_40_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_40_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_40_pat_count_3 <= _source_stream_conv2d_4_source_40_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_40_source_ram_renable <= 0;
        _stream_conv2d_4_source_40_idle <= 1;
      end 
      if((_stream_conv2d_4_source_40_source_pat_fsm_22 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_40_source_ram_renable <= 0;
        _stream_conv2d_4_source_40_idle <= 1;
      end 
      if(_set_flag_358) begin
        _stream_conv2d_4_source_41_source_mode <= 5'b10;
        _stream_conv2d_4_source_41_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_358) begin
        _source_stream_conv2d_4_source_41_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_41_pat_stride_0 <= 1;
      end 
      if(_set_flag_358) begin
        _source_stream_conv2d_4_source_41_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_41_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_358) begin
        _source_stream_conv2d_4_source_41_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_41_pat_stride_2 <= 0;
      end 
      if(_set_flag_358) begin
        _source_stream_conv2d_4_source_41_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_41_pat_stride_3 <= 0;
      end 
      if(_set_flag_358) begin
        _stream_conv2d_4_source_41_source_sel <= 24;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_41_source_offset_buf <= _stream_conv2d_4_source_41_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_count_0 <= _source_stream_conv2d_4_source_41_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_count_1 <= _source_stream_conv2d_4_source_41_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_count_2 <= _source_stream_conv2d_4_source_41_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_count_3 <= _source_stream_conv2d_4_source_41_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_size_buf_0 <= _source_stream_conv2d_4_source_41_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_size_buf_1 <= _source_stream_conv2d_4_source_41_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_size_buf_2 <= _source_stream_conv2d_4_source_41_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_size_buf_3 <= _source_stream_conv2d_4_source_41_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_stride_buf_0 <= _source_stream_conv2d_4_source_41_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_stride_buf_1 <= _source_stream_conv2d_4_source_41_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_stride_buf_2 <= _source_stream_conv2d_4_source_41_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_stride_buf_3 <= _source_stream_conv2d_4_source_41_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1340 <= _stream_conv2d_4_source_41_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_41_idle <= 0;
        _stream_conv2d_4_source_41_source_ram_raddr <= _stream_conv2d_4_source_41_source_pat_all_offset;
        _stream_conv2d_4_source_41_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_0 <= _source_stream_conv2d_4_source_41_pat_cur_offset_0 + _source_stream_conv2d_4_source_41_pat_stride_buf_0;
        _source_stream_conv2d_4_source_41_pat_count_0 <= _source_stream_conv2d_4_source_41_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && (_source_stream_conv2d_4_source_41_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_41_pat_count_0 <= _source_stream_conv2d_4_source_41_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && (_source_stream_conv2d_4_source_41_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_1 <= _source_stream_conv2d_4_source_41_pat_cur_offset_1 + _source_stream_conv2d_4_source_41_pat_stride_buf_1;
        _source_stream_conv2d_4_source_41_pat_count_1 <= _source_stream_conv2d_4_source_41_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && (_source_stream_conv2d_4_source_41_pat_count_0 == 0) && (_source_stream_conv2d_4_source_41_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_41_pat_count_1 <= _source_stream_conv2d_4_source_41_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && ((_source_stream_conv2d_4_source_41_pat_count_0 == 0) && (_source_stream_conv2d_4_source_41_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_2 <= _source_stream_conv2d_4_source_41_pat_cur_offset_2 + _source_stream_conv2d_4_source_41_pat_stride_buf_2;
        _source_stream_conv2d_4_source_41_pat_count_2 <= _source_stream_conv2d_4_source_41_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && ((_source_stream_conv2d_4_source_41_pat_count_0 == 0) && (_source_stream_conv2d_4_source_41_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_41_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_41_pat_count_2 <= _source_stream_conv2d_4_source_41_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && ((_source_stream_conv2d_4_source_41_pat_count_0 == 0) && (_source_stream_conv2d_4_source_41_pat_count_1 == 0) && (_source_stream_conv2d_4_source_41_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_3 <= _source_stream_conv2d_4_source_41_pat_cur_offset_3 + _source_stream_conv2d_4_source_41_pat_stride_buf_3;
        _source_stream_conv2d_4_source_41_pat_count_3 <= _source_stream_conv2d_4_source_41_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && ((_source_stream_conv2d_4_source_41_pat_count_0 == 0) && (_source_stream_conv2d_4_source_41_pat_count_1 == 0) && (_source_stream_conv2d_4_source_41_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_41_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_41_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_41_pat_count_3 <= _source_stream_conv2d_4_source_41_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_41_source_ram_renable <= 0;
        _stream_conv2d_4_source_41_idle <= 1;
      end 
      if((_stream_conv2d_4_source_41_source_pat_fsm_23 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_41_source_ram_renable <= 0;
        _stream_conv2d_4_source_41_idle <= 1;
      end 
      if(_set_flag_361) begin
        _stream_conv2d_4_source_42_source_mode <= 5'b10;
        _stream_conv2d_4_source_42_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_361) begin
        _source_stream_conv2d_4_source_42_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_42_pat_stride_0 <= 1;
      end 
      if(_set_flag_361) begin
        _source_stream_conv2d_4_source_42_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_42_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_361) begin
        _source_stream_conv2d_4_source_42_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_42_pat_stride_2 <= 0;
      end 
      if(_set_flag_361) begin
        _source_stream_conv2d_4_source_42_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_42_pat_stride_3 <= 0;
      end 
      if(_set_flag_361) begin
        _stream_conv2d_4_source_42_source_sel <= 25;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_42_source_offset_buf <= _stream_conv2d_4_source_42_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_count_0 <= _source_stream_conv2d_4_source_42_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_count_1 <= _source_stream_conv2d_4_source_42_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_count_2 <= _source_stream_conv2d_4_source_42_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_count_3 <= _source_stream_conv2d_4_source_42_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_size_buf_0 <= _source_stream_conv2d_4_source_42_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_size_buf_1 <= _source_stream_conv2d_4_source_42_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_size_buf_2 <= _source_stream_conv2d_4_source_42_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_size_buf_3 <= _source_stream_conv2d_4_source_42_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_stride_buf_0 <= _source_stream_conv2d_4_source_42_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_stride_buf_1 <= _source_stream_conv2d_4_source_42_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_stride_buf_2 <= _source_stream_conv2d_4_source_42_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_stride_buf_3 <= _source_stream_conv2d_4_source_42_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1341 <= _stream_conv2d_4_source_42_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_42_idle <= 0;
        _stream_conv2d_4_source_42_source_ram_raddr <= _stream_conv2d_4_source_42_source_pat_all_offset;
        _stream_conv2d_4_source_42_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_0 <= _source_stream_conv2d_4_source_42_pat_cur_offset_0 + _source_stream_conv2d_4_source_42_pat_stride_buf_0;
        _source_stream_conv2d_4_source_42_pat_count_0 <= _source_stream_conv2d_4_source_42_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && (_source_stream_conv2d_4_source_42_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_42_pat_count_0 <= _source_stream_conv2d_4_source_42_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && (_source_stream_conv2d_4_source_42_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_1 <= _source_stream_conv2d_4_source_42_pat_cur_offset_1 + _source_stream_conv2d_4_source_42_pat_stride_buf_1;
        _source_stream_conv2d_4_source_42_pat_count_1 <= _source_stream_conv2d_4_source_42_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && (_source_stream_conv2d_4_source_42_pat_count_0 == 0) && (_source_stream_conv2d_4_source_42_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_42_pat_count_1 <= _source_stream_conv2d_4_source_42_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && ((_source_stream_conv2d_4_source_42_pat_count_0 == 0) && (_source_stream_conv2d_4_source_42_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_2 <= _source_stream_conv2d_4_source_42_pat_cur_offset_2 + _source_stream_conv2d_4_source_42_pat_stride_buf_2;
        _source_stream_conv2d_4_source_42_pat_count_2 <= _source_stream_conv2d_4_source_42_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && ((_source_stream_conv2d_4_source_42_pat_count_0 == 0) && (_source_stream_conv2d_4_source_42_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_42_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_42_pat_count_2 <= _source_stream_conv2d_4_source_42_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && ((_source_stream_conv2d_4_source_42_pat_count_0 == 0) && (_source_stream_conv2d_4_source_42_pat_count_1 == 0) && (_source_stream_conv2d_4_source_42_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_3 <= _source_stream_conv2d_4_source_42_pat_cur_offset_3 + _source_stream_conv2d_4_source_42_pat_stride_buf_3;
        _source_stream_conv2d_4_source_42_pat_count_3 <= _source_stream_conv2d_4_source_42_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && ((_source_stream_conv2d_4_source_42_pat_count_0 == 0) && (_source_stream_conv2d_4_source_42_pat_count_1 == 0) && (_source_stream_conv2d_4_source_42_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_42_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_42_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_42_pat_count_3 <= _source_stream_conv2d_4_source_42_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_42_source_ram_renable <= 0;
        _stream_conv2d_4_source_42_idle <= 1;
      end 
      if((_stream_conv2d_4_source_42_source_pat_fsm_24 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_42_source_ram_renable <= 0;
        _stream_conv2d_4_source_42_idle <= 1;
      end 
      if(_set_flag_364) begin
        _stream_conv2d_4_source_43_source_mode <= 5'b10;
        _stream_conv2d_4_source_43_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_364) begin
        _source_stream_conv2d_4_source_43_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_43_pat_stride_0 <= 1;
      end 
      if(_set_flag_364) begin
        _source_stream_conv2d_4_source_43_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_43_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_364) begin
        _source_stream_conv2d_4_source_43_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_43_pat_stride_2 <= 0;
      end 
      if(_set_flag_364) begin
        _source_stream_conv2d_4_source_43_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_43_pat_stride_3 <= 0;
      end 
      if(_set_flag_364) begin
        _stream_conv2d_4_source_43_source_sel <= 26;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_43_source_offset_buf <= _stream_conv2d_4_source_43_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_count_0 <= _source_stream_conv2d_4_source_43_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_count_1 <= _source_stream_conv2d_4_source_43_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_count_2 <= _source_stream_conv2d_4_source_43_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_count_3 <= _source_stream_conv2d_4_source_43_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_size_buf_0 <= _source_stream_conv2d_4_source_43_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_size_buf_1 <= _source_stream_conv2d_4_source_43_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_size_buf_2 <= _source_stream_conv2d_4_source_43_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_size_buf_3 <= _source_stream_conv2d_4_source_43_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_stride_buf_0 <= _source_stream_conv2d_4_source_43_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_stride_buf_1 <= _source_stream_conv2d_4_source_43_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_stride_buf_2 <= _source_stream_conv2d_4_source_43_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_stride_buf_3 <= _source_stream_conv2d_4_source_43_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1342 <= _stream_conv2d_4_source_43_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_43_idle <= 0;
        _stream_conv2d_4_source_43_source_ram_raddr <= _stream_conv2d_4_source_43_source_pat_all_offset;
        _stream_conv2d_4_source_43_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_0 <= _source_stream_conv2d_4_source_43_pat_cur_offset_0 + _source_stream_conv2d_4_source_43_pat_stride_buf_0;
        _source_stream_conv2d_4_source_43_pat_count_0 <= _source_stream_conv2d_4_source_43_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && (_source_stream_conv2d_4_source_43_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_43_pat_count_0 <= _source_stream_conv2d_4_source_43_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && (_source_stream_conv2d_4_source_43_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_1 <= _source_stream_conv2d_4_source_43_pat_cur_offset_1 + _source_stream_conv2d_4_source_43_pat_stride_buf_1;
        _source_stream_conv2d_4_source_43_pat_count_1 <= _source_stream_conv2d_4_source_43_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && (_source_stream_conv2d_4_source_43_pat_count_0 == 0) && (_source_stream_conv2d_4_source_43_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_43_pat_count_1 <= _source_stream_conv2d_4_source_43_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && ((_source_stream_conv2d_4_source_43_pat_count_0 == 0) && (_source_stream_conv2d_4_source_43_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_2 <= _source_stream_conv2d_4_source_43_pat_cur_offset_2 + _source_stream_conv2d_4_source_43_pat_stride_buf_2;
        _source_stream_conv2d_4_source_43_pat_count_2 <= _source_stream_conv2d_4_source_43_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && ((_source_stream_conv2d_4_source_43_pat_count_0 == 0) && (_source_stream_conv2d_4_source_43_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_43_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_43_pat_count_2 <= _source_stream_conv2d_4_source_43_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && ((_source_stream_conv2d_4_source_43_pat_count_0 == 0) && (_source_stream_conv2d_4_source_43_pat_count_1 == 0) && (_source_stream_conv2d_4_source_43_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_3 <= _source_stream_conv2d_4_source_43_pat_cur_offset_3 + _source_stream_conv2d_4_source_43_pat_stride_buf_3;
        _source_stream_conv2d_4_source_43_pat_count_3 <= _source_stream_conv2d_4_source_43_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && ((_source_stream_conv2d_4_source_43_pat_count_0 == 0) && (_source_stream_conv2d_4_source_43_pat_count_1 == 0) && (_source_stream_conv2d_4_source_43_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_43_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_43_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_43_pat_count_3 <= _source_stream_conv2d_4_source_43_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_43_source_ram_renable <= 0;
        _stream_conv2d_4_source_43_idle <= 1;
      end 
      if((_stream_conv2d_4_source_43_source_pat_fsm_25 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_43_source_ram_renable <= 0;
        _stream_conv2d_4_source_43_idle <= 1;
      end 
      if(_set_flag_367) begin
        _stream_conv2d_4_source_44_source_mode <= 5'b10;
        _stream_conv2d_4_source_44_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_367) begin
        _source_stream_conv2d_4_source_44_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_44_pat_stride_0 <= 1;
      end 
      if(_set_flag_367) begin
        _source_stream_conv2d_4_source_44_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_44_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_367) begin
        _source_stream_conv2d_4_source_44_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_44_pat_stride_2 <= 0;
      end 
      if(_set_flag_367) begin
        _source_stream_conv2d_4_source_44_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_44_pat_stride_3 <= 0;
      end 
      if(_set_flag_367) begin
        _stream_conv2d_4_source_44_source_sel <= 27;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_44_source_offset_buf <= _stream_conv2d_4_source_44_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_count_0 <= _source_stream_conv2d_4_source_44_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_count_1 <= _source_stream_conv2d_4_source_44_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_count_2 <= _source_stream_conv2d_4_source_44_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_count_3 <= _source_stream_conv2d_4_source_44_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_size_buf_0 <= _source_stream_conv2d_4_source_44_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_size_buf_1 <= _source_stream_conv2d_4_source_44_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_size_buf_2 <= _source_stream_conv2d_4_source_44_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_size_buf_3 <= _source_stream_conv2d_4_source_44_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_stride_buf_0 <= _source_stream_conv2d_4_source_44_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_stride_buf_1 <= _source_stream_conv2d_4_source_44_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_stride_buf_2 <= _source_stream_conv2d_4_source_44_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_stride_buf_3 <= _source_stream_conv2d_4_source_44_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1343 <= _stream_conv2d_4_source_44_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_44_idle <= 0;
        _stream_conv2d_4_source_44_source_ram_raddr <= _stream_conv2d_4_source_44_source_pat_all_offset;
        _stream_conv2d_4_source_44_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_0 <= _source_stream_conv2d_4_source_44_pat_cur_offset_0 + _source_stream_conv2d_4_source_44_pat_stride_buf_0;
        _source_stream_conv2d_4_source_44_pat_count_0 <= _source_stream_conv2d_4_source_44_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && (_source_stream_conv2d_4_source_44_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_44_pat_count_0 <= _source_stream_conv2d_4_source_44_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && (_source_stream_conv2d_4_source_44_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_1 <= _source_stream_conv2d_4_source_44_pat_cur_offset_1 + _source_stream_conv2d_4_source_44_pat_stride_buf_1;
        _source_stream_conv2d_4_source_44_pat_count_1 <= _source_stream_conv2d_4_source_44_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && (_source_stream_conv2d_4_source_44_pat_count_0 == 0) && (_source_stream_conv2d_4_source_44_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_44_pat_count_1 <= _source_stream_conv2d_4_source_44_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && ((_source_stream_conv2d_4_source_44_pat_count_0 == 0) && (_source_stream_conv2d_4_source_44_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_2 <= _source_stream_conv2d_4_source_44_pat_cur_offset_2 + _source_stream_conv2d_4_source_44_pat_stride_buf_2;
        _source_stream_conv2d_4_source_44_pat_count_2 <= _source_stream_conv2d_4_source_44_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && ((_source_stream_conv2d_4_source_44_pat_count_0 == 0) && (_source_stream_conv2d_4_source_44_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_44_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_44_pat_count_2 <= _source_stream_conv2d_4_source_44_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && ((_source_stream_conv2d_4_source_44_pat_count_0 == 0) && (_source_stream_conv2d_4_source_44_pat_count_1 == 0) && (_source_stream_conv2d_4_source_44_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_3 <= _source_stream_conv2d_4_source_44_pat_cur_offset_3 + _source_stream_conv2d_4_source_44_pat_stride_buf_3;
        _source_stream_conv2d_4_source_44_pat_count_3 <= _source_stream_conv2d_4_source_44_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && ((_source_stream_conv2d_4_source_44_pat_count_0 == 0) && (_source_stream_conv2d_4_source_44_pat_count_1 == 0) && (_source_stream_conv2d_4_source_44_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_44_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_44_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_44_pat_count_3 <= _source_stream_conv2d_4_source_44_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_44_source_ram_renable <= 0;
        _stream_conv2d_4_source_44_idle <= 1;
      end 
      if((_stream_conv2d_4_source_44_source_pat_fsm_26 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_44_source_ram_renable <= 0;
        _stream_conv2d_4_source_44_idle <= 1;
      end 
      if(_set_flag_370) begin
        _stream_conv2d_4_source_45_source_mode <= 5'b10;
        _stream_conv2d_4_source_45_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_370) begin
        _source_stream_conv2d_4_source_45_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_45_pat_stride_0 <= 1;
      end 
      if(_set_flag_370) begin
        _source_stream_conv2d_4_source_45_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_45_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_370) begin
        _source_stream_conv2d_4_source_45_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_45_pat_stride_2 <= 0;
      end 
      if(_set_flag_370) begin
        _source_stream_conv2d_4_source_45_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_45_pat_stride_3 <= 0;
      end 
      if(_set_flag_370) begin
        _stream_conv2d_4_source_45_source_sel <= 28;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_45_source_offset_buf <= _stream_conv2d_4_source_45_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_count_0 <= _source_stream_conv2d_4_source_45_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_count_1 <= _source_stream_conv2d_4_source_45_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_count_2 <= _source_stream_conv2d_4_source_45_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_count_3 <= _source_stream_conv2d_4_source_45_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_size_buf_0 <= _source_stream_conv2d_4_source_45_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_size_buf_1 <= _source_stream_conv2d_4_source_45_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_size_buf_2 <= _source_stream_conv2d_4_source_45_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_size_buf_3 <= _source_stream_conv2d_4_source_45_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_stride_buf_0 <= _source_stream_conv2d_4_source_45_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_stride_buf_1 <= _source_stream_conv2d_4_source_45_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_stride_buf_2 <= _source_stream_conv2d_4_source_45_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_stride_buf_3 <= _source_stream_conv2d_4_source_45_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1344 <= _stream_conv2d_4_source_45_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_45_idle <= 0;
        _stream_conv2d_4_source_45_source_ram_raddr <= _stream_conv2d_4_source_45_source_pat_all_offset;
        _stream_conv2d_4_source_45_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_0 <= _source_stream_conv2d_4_source_45_pat_cur_offset_0 + _source_stream_conv2d_4_source_45_pat_stride_buf_0;
        _source_stream_conv2d_4_source_45_pat_count_0 <= _source_stream_conv2d_4_source_45_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && (_source_stream_conv2d_4_source_45_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_45_pat_count_0 <= _source_stream_conv2d_4_source_45_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && (_source_stream_conv2d_4_source_45_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_1 <= _source_stream_conv2d_4_source_45_pat_cur_offset_1 + _source_stream_conv2d_4_source_45_pat_stride_buf_1;
        _source_stream_conv2d_4_source_45_pat_count_1 <= _source_stream_conv2d_4_source_45_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && (_source_stream_conv2d_4_source_45_pat_count_0 == 0) && (_source_stream_conv2d_4_source_45_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_45_pat_count_1 <= _source_stream_conv2d_4_source_45_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && ((_source_stream_conv2d_4_source_45_pat_count_0 == 0) && (_source_stream_conv2d_4_source_45_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_2 <= _source_stream_conv2d_4_source_45_pat_cur_offset_2 + _source_stream_conv2d_4_source_45_pat_stride_buf_2;
        _source_stream_conv2d_4_source_45_pat_count_2 <= _source_stream_conv2d_4_source_45_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && ((_source_stream_conv2d_4_source_45_pat_count_0 == 0) && (_source_stream_conv2d_4_source_45_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_45_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_45_pat_count_2 <= _source_stream_conv2d_4_source_45_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && ((_source_stream_conv2d_4_source_45_pat_count_0 == 0) && (_source_stream_conv2d_4_source_45_pat_count_1 == 0) && (_source_stream_conv2d_4_source_45_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_3 <= _source_stream_conv2d_4_source_45_pat_cur_offset_3 + _source_stream_conv2d_4_source_45_pat_stride_buf_3;
        _source_stream_conv2d_4_source_45_pat_count_3 <= _source_stream_conv2d_4_source_45_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && ((_source_stream_conv2d_4_source_45_pat_count_0 == 0) && (_source_stream_conv2d_4_source_45_pat_count_1 == 0) && (_source_stream_conv2d_4_source_45_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_45_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_45_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_45_pat_count_3 <= _source_stream_conv2d_4_source_45_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_45_source_ram_renable <= 0;
        _stream_conv2d_4_source_45_idle <= 1;
      end 
      if((_stream_conv2d_4_source_45_source_pat_fsm_27 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_45_source_ram_renable <= 0;
        _stream_conv2d_4_source_45_idle <= 1;
      end 
      if(_set_flag_373) begin
        _stream_conv2d_4_source_46_source_mode <= 5'b10;
        _stream_conv2d_4_source_46_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_373) begin
        _source_stream_conv2d_4_source_46_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_46_pat_stride_0 <= 1;
      end 
      if(_set_flag_373) begin
        _source_stream_conv2d_4_source_46_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_46_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_373) begin
        _source_stream_conv2d_4_source_46_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_46_pat_stride_2 <= 0;
      end 
      if(_set_flag_373) begin
        _source_stream_conv2d_4_source_46_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_46_pat_stride_3 <= 0;
      end 
      if(_set_flag_373) begin
        _stream_conv2d_4_source_46_source_sel <= 29;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_46_source_offset_buf <= _stream_conv2d_4_source_46_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_count_0 <= _source_stream_conv2d_4_source_46_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_count_1 <= _source_stream_conv2d_4_source_46_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_count_2 <= _source_stream_conv2d_4_source_46_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_count_3 <= _source_stream_conv2d_4_source_46_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_size_buf_0 <= _source_stream_conv2d_4_source_46_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_size_buf_1 <= _source_stream_conv2d_4_source_46_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_size_buf_2 <= _source_stream_conv2d_4_source_46_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_size_buf_3 <= _source_stream_conv2d_4_source_46_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_stride_buf_0 <= _source_stream_conv2d_4_source_46_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_stride_buf_1 <= _source_stream_conv2d_4_source_46_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_stride_buf_2 <= _source_stream_conv2d_4_source_46_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_stride_buf_3 <= _source_stream_conv2d_4_source_46_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1345 <= _stream_conv2d_4_source_46_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_46_idle <= 0;
        _stream_conv2d_4_source_46_source_ram_raddr <= _stream_conv2d_4_source_46_source_pat_all_offset;
        _stream_conv2d_4_source_46_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_0 <= _source_stream_conv2d_4_source_46_pat_cur_offset_0 + _source_stream_conv2d_4_source_46_pat_stride_buf_0;
        _source_stream_conv2d_4_source_46_pat_count_0 <= _source_stream_conv2d_4_source_46_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && (_source_stream_conv2d_4_source_46_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_46_pat_count_0 <= _source_stream_conv2d_4_source_46_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && (_source_stream_conv2d_4_source_46_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_1 <= _source_stream_conv2d_4_source_46_pat_cur_offset_1 + _source_stream_conv2d_4_source_46_pat_stride_buf_1;
        _source_stream_conv2d_4_source_46_pat_count_1 <= _source_stream_conv2d_4_source_46_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && (_source_stream_conv2d_4_source_46_pat_count_0 == 0) && (_source_stream_conv2d_4_source_46_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_46_pat_count_1 <= _source_stream_conv2d_4_source_46_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && ((_source_stream_conv2d_4_source_46_pat_count_0 == 0) && (_source_stream_conv2d_4_source_46_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_2 <= _source_stream_conv2d_4_source_46_pat_cur_offset_2 + _source_stream_conv2d_4_source_46_pat_stride_buf_2;
        _source_stream_conv2d_4_source_46_pat_count_2 <= _source_stream_conv2d_4_source_46_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && ((_source_stream_conv2d_4_source_46_pat_count_0 == 0) && (_source_stream_conv2d_4_source_46_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_46_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_46_pat_count_2 <= _source_stream_conv2d_4_source_46_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && ((_source_stream_conv2d_4_source_46_pat_count_0 == 0) && (_source_stream_conv2d_4_source_46_pat_count_1 == 0) && (_source_stream_conv2d_4_source_46_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_3 <= _source_stream_conv2d_4_source_46_pat_cur_offset_3 + _source_stream_conv2d_4_source_46_pat_stride_buf_3;
        _source_stream_conv2d_4_source_46_pat_count_3 <= _source_stream_conv2d_4_source_46_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && ((_source_stream_conv2d_4_source_46_pat_count_0 == 0) && (_source_stream_conv2d_4_source_46_pat_count_1 == 0) && (_source_stream_conv2d_4_source_46_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_46_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_46_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_46_pat_count_3 <= _source_stream_conv2d_4_source_46_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_46_source_ram_renable <= 0;
        _stream_conv2d_4_source_46_idle <= 1;
      end 
      if((_stream_conv2d_4_source_46_source_pat_fsm_28 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_46_source_ram_renable <= 0;
        _stream_conv2d_4_source_46_idle <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_377 <= _set_flag_376;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_378 <= _tmp_377;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_379 <= _tmp_378;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_380 <= _tmp_379;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_381 <= _tmp_380;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_382 <= _tmp_381;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_383 <= _tmp_382;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_384 <= _tmp_383;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_385 <= _tmp_384;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_386 <= _tmp_385;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_387 <= _tmp_386;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_388 <= _tmp_387;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_389 <= _tmp_388;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_390 <= _tmp_389;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_391 <= _tmp_390;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_392 <= _tmp_391;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_393 <= _tmp_392;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_394 <= _tmp_393;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_395 <= _tmp_394;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_396 <= _tmp_395;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_397 <= _tmp_396;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_398 <= _tmp_397;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_399 <= _tmp_398;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_400 <= _tmp_399;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_401 <= _tmp_400;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_402 <= _tmp_401;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_403 <= _tmp_402;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_404 <= _tmp_403;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_405 <= _tmp_404;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_406 <= _tmp_405;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_407 <= _tmp_406;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_408 <= _tmp_407;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_409 <= _tmp_408;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_410 <= _tmp_409;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_411 <= _tmp_410;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_412 <= _tmp_411;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_415 <= _tmp_414;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_416 <= _tmp_415;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_417 <= _tmp_416;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_418 <= _tmp_417;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_419 <= _tmp_418;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_420 <= _tmp_419;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_421 <= _tmp_420;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_422 <= _tmp_421;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_423 <= _tmp_422;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_424 <= _tmp_423;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_425 <= _tmp_424;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_426 <= _tmp_425;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_427 <= _tmp_426;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_428 <= _tmp_427;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_429 <= _tmp_428;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_430 <= _tmp_429;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_431 <= _tmp_430;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_432 <= _tmp_431;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_433 <= _tmp_432;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_434 <= _tmp_433;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_435 <= _tmp_434;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_436 <= _tmp_435;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_437 <= _tmp_436;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_438 <= _tmp_437;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_439 <= _tmp_438;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_440 <= _tmp_439;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_441 <= _tmp_440;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_442 <= _tmp_441;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_443 <= _tmp_442;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_444 <= _tmp_443;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_445 <= _tmp_444;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_446 <= _tmp_445;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_447 <= _tmp_446;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_448 <= _tmp_447;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_449 <= _tmp_448;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_450 <= _tmp_449;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_451 <= conv2d_4_next_stream_num_ops;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_452 <= _tmp_451;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_453 <= _tmp_452;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_454 <= _tmp_453;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_455 <= _tmp_454;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_456 <= _tmp_455;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_457 <= _tmp_456;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_458 <= _tmp_457;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_459 <= _tmp_458;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_460 <= _tmp_459;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_461 <= _tmp_460;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_462 <= _tmp_461;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_463 <= _tmp_462;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_464 <= _tmp_463;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_465 <= _tmp_464;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_466 <= _tmp_465;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_467 <= _tmp_466;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_468 <= _tmp_467;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_469 <= _tmp_468;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_470 <= _tmp_469;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_471 <= _tmp_470;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_472 <= _tmp_471;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_473 <= _tmp_472;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_474 <= _tmp_473;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_475 <= _tmp_474;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_476 <= _tmp_475;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_477 <= _tmp_476;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_478 <= _tmp_477;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_479 <= _tmp_478;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_480 <= _tmp_479;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_481 <= _tmp_480;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_482 <= _tmp_481;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_483 <= _tmp_482;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_484 <= _tmp_483;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_485 <= _tmp_484;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_486 <= _tmp_485;
      end 
      if(_tmp_412) begin
        _stream_conv2d_4_sink_89_sink_mode <= 5'b1;
        _stream_conv2d_4_sink_89_sink_offset <= _tmp_450;
        _stream_conv2d_4_sink_89_sink_size <= _tmp_486;
        _stream_conv2d_4_sink_89_sink_stride <= 1;
      end 
      if(_tmp_412) begin
        _stream_conv2d_4_sink_89_sink_sel <= 30;
      end 
      if(_stream_conv2d_4_sink_start && _stream_conv2d_4_sink_89_sink_mode & 5'b1 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_89_sink_offset_buf <= _stream_conv2d_4_sink_89_sink_offset;
        _stream_conv2d_4_sink_89_sink_size_buf <= _stream_conv2d_4_sink_89_sink_size;
        _stream_conv2d_4_sink_89_sink_stride_buf <= _stream_conv2d_4_sink_89_sink_stride;
      end 
      if((_stream_conv2d_4_sink_89_sink_fsm_29 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_89_sink_waddr <= _stream_conv2d_4_sink_89_sink_offset_buf - _stream_conv2d_4_sink_89_sink_stride_buf;
        _stream_conv2d_4_sink_89_sink_count <= _stream_conv2d_4_sink_89_sink_size_buf;
      end 
      if((_stream_conv2d_4_sink_89_sink_fsm_29 == 2) && stream_conv2d_4_sink_90_data && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_89_sink_waddr <= _stream_conv2d_4_sink_89_sink_waddr + _stream_conv2d_4_sink_89_sink_stride_buf;
        _stream_conv2d_4_sink_89_sink_wdata <= stream_conv2d_4_sink_89_data;
        _stream_conv2d_4_sink_89_sink_wenable <= 1;
        _stream_conv2d_4_sink_89_sink_count <= _stream_conv2d_4_sink_89_sink_count - 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1882 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1883 <= _tmp_1882;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1884 <= _tmp_1883;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1885 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1886 <= _tmp_1885;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1887 <= _tmp_1886;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1887) begin
        __variable_wdata_951 <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1888 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1889 <= _tmp_1888;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1890 <= _tmp_1889;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1891 <= _tmp_1890;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1891) begin
        __variable_wdata_951 <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1894 <= _tmp_1893;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1897 <= _tmp_1896;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1897) begin
        __variable_wdata_951 <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1898 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1899 <= _tmp_1898;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1900 <= _tmp_1899;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1901 <= _tmp_1900;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1902 <= _tmp_1901;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1903 <= _tmp_1902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1904 <= _tmp_1903;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1905 <= _tmp_1904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1906 <= _tmp_1905;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1907 <= _tmp_1906;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1908 <= _tmp_1907;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1909 <= _tmp_1908;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1910 <= _tmp_1909;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1911 <= _tmp_1910;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1912 <= _tmp_1911;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1913 <= _tmp_1912;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1914 <= _tmp_1913;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1915 <= _tmp_1914;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1916 <= _tmp_1915;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1917 <= _tmp_1916;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1918 <= _tmp_1917;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1919 <= _tmp_1918;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1920 <= _tmp_1919;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1921 <= _tmp_1920;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1922 <= _tmp_1921;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1923 <= _tmp_1922;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1924 <= _tmp_1923;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1925 <= _tmp_1924;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1926 <= _tmp_1925;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1927 <= _tmp_1926;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1928 <= _tmp_1927;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1929 <= _tmp_1928;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1930 <= _tmp_1929;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1931 <= _tmp_1930;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1932 <= _tmp_1931;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1933 <= _tmp_1932;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1934 <= _stream_conv2d_4_source_stop;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1935 <= _tmp_1934;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1936 <= _tmp_1935;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1937 <= _tmp_1936;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1938 <= _tmp_1937;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1939 <= _tmp_1938;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1940 <= _tmp_1939;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1941 <= _tmp_1940;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1942 <= _tmp_1941;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1943 <= _tmp_1942;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1944 <= _tmp_1943;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1945 <= _tmp_1944;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1946 <= _tmp_1945;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1947 <= _tmp_1946;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1948 <= _tmp_1947;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1949 <= _tmp_1948;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1950 <= _tmp_1949;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1951 <= _tmp_1950;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1952 <= _tmp_1951;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1953 <= _tmp_1952;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1954 <= _tmp_1953;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1955 <= _tmp_1954;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1956 <= _tmp_1955;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1957 <= _tmp_1956;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1958 <= _tmp_1957;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1959 <= _tmp_1958;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1960 <= _tmp_1959;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1961 <= _tmp_1960;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1962 <= _tmp_1961;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1963 <= _tmp_1962;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1964 <= _tmp_1963;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1965 <= _tmp_1964;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1966 <= _tmp_1965;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1967 <= _tmp_1966;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1968 <= _tmp_1967;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1969 <= _tmp_1968;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1970 <= _stream_conv2d_4_source_busy;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1971 <= _tmp_1970;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1972 <= _tmp_1971;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1973 <= _tmp_1972;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1974 <= _tmp_1973;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1975 <= _tmp_1974;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1976 <= _tmp_1975;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1977 <= _tmp_1976;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1978 <= _tmp_1977;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1979 <= _tmp_1978;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1980 <= _tmp_1979;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1981 <= _tmp_1980;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1982 <= _tmp_1981;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1983 <= _tmp_1982;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1984 <= _tmp_1983;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1985 <= _tmp_1984;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1986 <= _tmp_1985;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1987 <= _tmp_1986;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1988 <= _tmp_1987;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1989 <= _tmp_1988;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1990 <= _tmp_1989;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1991 <= _tmp_1990;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1992 <= _tmp_1991;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1993 <= _tmp_1992;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1994 <= _tmp_1993;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1995 <= _tmp_1994;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1996 <= _tmp_1995;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1997 <= _tmp_1996;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1998 <= _tmp_1997;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1999 <= _tmp_1998;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_2000 <= _tmp_1999;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_2001 <= _tmp_2000;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_2002 <= _tmp_2001;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_2003 <= _tmp_2002;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_2004 <= _tmp_2003;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_2005 <= _tmp_2004;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_2006 <= _stream_conv2d_4_sink_busy;
      end 
      if(!_stream_conv2d_4_sink_busy && _tmp_2006) begin
        _stream_conv2d_4_busy_reg <= 0;
      end 
      if(_stream_conv2d_4_source_busy) begin
        _stream_conv2d_4_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_conv2d_4_fsm_1 = 1;
  localparam _stream_conv2d_4_fsm_2 = 2;
  localparam _stream_conv2d_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_init;
      _stream_conv2d_4_source_start <= 0;
      _stream_conv2d_4_source_busy <= 0;
      _stream_conv2d_4_stream_ivalid <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _tmp_1884) begin
        _stream_conv2d_4_stream_ivalid <= 1;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1894) begin
        _stream_conv2d_4_stream_ivalid <= 0;
      end 
      case(_stream_conv2d_4_fsm)
        _stream_conv2d_4_fsm_init: begin
          if(_stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_source_start <= 1;
          end 
          if(_stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_1;
          end 
        end
        _stream_conv2d_4_fsm_1: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_start <= 0;
            _stream_conv2d_4_source_busy <= 1;
          end 
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_2;
          end 
        end
        _stream_conv2d_4_fsm_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_3;
          end 
        end
        _stream_conv2d_4_fsm_3: begin
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_38_idle && _stream_conv2d_4_source_39_idle && _stream_conv2d_4_source_40_idle && _stream_conv2d_4_source_41_idle && _stream_conv2d_4_source_42_idle && _stream_conv2d_4_source_43_idle && _stream_conv2d_4_source_44_idle && _stream_conv2d_4_source_45_idle && _stream_conv2d_4_source_46_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3))) begin
            _stream_conv2d_4_source_busy <= 0;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_38_idle && _stream_conv2d_4_source_39_idle && _stream_conv2d_4_source_40_idle && _stream_conv2d_4_source_41_idle && _stream_conv2d_4_source_42_idle && _stream_conv2d_4_source_43_idle && _stream_conv2d_4_source_44_idle && _stream_conv2d_4_source_45_idle && _stream_conv2d_4_source_46_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3)) && _stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_source_start <= 1;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_38_idle && _stream_conv2d_4_source_39_idle && _stream_conv2d_4_source_40_idle && _stream_conv2d_4_source_41_idle && _stream_conv2d_4_source_42_idle && _stream_conv2d_4_source_43_idle && _stream_conv2d_4_source_44_idle && _stream_conv2d_4_source_45_idle && _stream_conv2d_4_source_46_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3))) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_init;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_38_idle && _stream_conv2d_4_source_39_idle && _stream_conv2d_4_source_40_idle && _stream_conv2d_4_source_41_idle && _stream_conv2d_4_source_42_idle && _stream_conv2d_4_source_43_idle && _stream_conv2d_4_source_44_idle && _stream_conv2d_4_source_45_idle && _stream_conv2d_4_source_46_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3)) && _stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
      _stream_max_pool_serial_6_source_1_source_fifo_deq <= 0;
      _stream_max_pool_serial_6_source_1_idle <= 1;
      _stream_max_pool_serial_6_sink_6_sink_wenable <= 0;
      _stream_max_pool_serial_6_sink_6_sink_fifo_enq <= 0;
      _stream_max_pool_serial_6_sink_7_sink_wenable <= 0;
      _stream_max_pool_serial_6_sink_7_sink_fifo_enq <= 0;
      __stream_max_pool_serial_6_stream_ivalid_1 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_2 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_3 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_4 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_5 <= 0;
      _counter_data_2421 <= 1'sd0;
      _counter_count_2421 <= 1'sd0;
      __delay_data_3108__variable_2419 <= 0;
      __delay_data_3109_reinterpretcast_2428 <= 0;
      __delay_data_3111__variable_2420 <= 0;
      __delay_data_3114__variable_2417 <= 0;
      __delay_data_3117_reinterpretcast_2432 <= 0;
      _pointer_data_2424 <= 0;
      __delay_data_3110__delay_3109_reinterpretcast_2428 <= 0;
      __delay_data_3112__delay_3111__variable_2420 <= 0;
      __delay_data_3115__delay_3114__variable_2417 <= 0;
      __delay_data_3118__delay_3117_reinterpretcast_2432 <= 0;
      _cond_data_2434 <= 0;
      _cond_data_2439 <= 0;
      __delay_data_3113__delay_3112__delay_3111__variable_2420 <= 0;
      __delay_data_3116__delay_3115__delay_3114__variable_2417 <= 0;
      _stream_max_pool_serial_6_parameter_0_next_parameter_data <= 0;
      __variable_wdata_2417 <= 0;
      _stream_max_pool_serial_6_parameter_2_next_parameter_data <= 0;
      __variable_wdata_2419 <= 0;
      _stream_max_pool_serial_6_source_1_source_mode <= 5'b0;
      _stream_max_pool_serial_6_source_1_source_offset <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_3 <= 0;
      _stream_max_pool_serial_6_source_1_source_sel <= 0;
      _stream_max_pool_serial_6_source_1_source_offset_buf <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3 <= 0;
      __variable_wdata_2418 <= 0;
      _stream_max_pool_serial_6_source_1_source_ram_raddr <= 0;
      _tmp_2059 <= 0;
      _tmp_2060 <= 0;
      _tmp_2061 <= 0;
      _tmp_2062 <= 0;
      _tmp_2063 <= 0;
      _tmp_2064 <= 0;
      _tmp_2065 <= 0;
      _tmp_2068 <= 0;
      _tmp_2069 <= 0;
      _tmp_2070 <= 0;
      _tmp_2071 <= 0;
      _tmp_2072 <= 0;
      _tmp_2073 <= 0;
      _tmp_2074 <= 0;
      _tmp_2075 <= 0;
      _tmp_2076 <= 0;
      _tmp_2077 <= 0;
      _tmp_2078 <= 0;
      _tmp_2079 <= 0;
      _tmp_2080 <= 0;
      _tmp_2081 <= 0;
      _stream_max_pool_serial_6_sink_6_sink_mode <= 5'b0;
      _stream_max_pool_serial_6_sink_6_sink_offset <= 0;
      _stream_max_pool_serial_6_sink_6_sink_size <= 0;
      _stream_max_pool_serial_6_sink_6_sink_stride <= 0;
      _stream_max_pool_serial_6_sink_6_sink_sel <= 0;
      _stream_max_pool_serial_6_sink_6_sink_offset_buf <= 0;
      _stream_max_pool_serial_6_sink_6_sink_size_buf <= 0;
      _stream_max_pool_serial_6_sink_6_sink_stride_buf <= 0;
      _stream_max_pool_serial_6_sink_6_sink_waddr <= 0;
      _stream_max_pool_serial_6_sink_6_sink_count <= 0;
      _stream_max_pool_serial_6_sink_6_sink_wdata <= 0;
      _tmp_2123 <= 0;
      _tmp_2124 <= 0;
      _tmp_2125 <= 0;
      _tmp_2126 <= 0;
      _tmp_2127 <= 0;
      _tmp_2128 <= 0;
      __variable_wdata_2420 <= 0;
      _tmp_2129 <= 0;
      _tmp_2130 <= 0;
      _tmp_2131 <= 0;
      _tmp_2132 <= 0;
      _tmp_2135 <= 0;
      _tmp_2138 <= 0;
      _tmp_2139 <= 0;
      _tmp_2140 <= 0;
      _tmp_2141 <= 0;
      _tmp_2142 <= 0;
      _tmp_2143 <= 0;
      _tmp_2144 <= 0;
      _tmp_2145 <= 0;
      _tmp_2146 <= 0;
      _tmp_2147 <= 0;
      _tmp_2148 <= 0;
      _tmp_2149 <= 0;
      _tmp_2150 <= 0;
      _tmp_2151 <= 0;
      _tmp_2152 <= 0;
      _tmp_2153 <= 0;
      _tmp_2154 <= 0;
      _tmp_2155 <= 0;
      _tmp_2156 <= 0;
      _tmp_2157 <= 0;
      _tmp_2158 <= 0;
      _tmp_2159 <= 0;
      _tmp_2160 <= 0;
      _stream_max_pool_serial_6_busy_reg <= 0;
    end else begin
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_source_fifo_deq <= 0;
      end 
      _stream_max_pool_serial_6_source_1_idle <= _stream_max_pool_serial_6_source_1_idle;
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_wenable <= 0;
        _stream_max_pool_serial_6_sink_6_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_7_sink_wenable <= 0;
        _stream_max_pool_serial_6_sink_7_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_1 <= _stream_max_pool_serial_6_stream_ivalid;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_2 <= __stream_max_pool_serial_6_stream_ivalid_1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_3 <= __stream_max_pool_serial_6_stream_ivalid_2;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_4 <= __stream_max_pool_serial_6_stream_ivalid_3;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_5 <= __stream_max_pool_serial_6_stream_ivalid_4;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready && _counter_reset_cond_2421) begin
        _counter_data_2421 <= 1'sd0;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready) begin
        _counter_data_2421 <= _counter_current_count_2421;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready) begin
        _counter_count_2421 <= (_counter_current_count_2421 >= stream_max_pool_serial_6_parameter_0_data - 2'sd1)? _counter_current_count_2421 + 2'sd1 - stream_max_pool_serial_6_parameter_0_data : _counter_current_count_2421 + 2'sd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3108__variable_2419 <= stream_max_pool_serial_6_parameter_2_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3109_reinterpretcast_2428 <= _reinterpretcast_data_2428;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3111__variable_2420 <= stream_max_pool_serial_6__reduce_reset_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3114__variable_2417 <= stream_max_pool_serial_6_parameter_0_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3117_reinterpretcast_2432 <= _reinterpretcast_data_2432;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _pointer_data_2424 <= __delay_data_3108__variable_2419[_counter_data_2421];
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3110__delay_3109_reinterpretcast_2428 <= __delay_data_3109_reinterpretcast_2428;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3112__delay_3111__variable_2420 <= __delay_data_3111__variable_2420;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3115__delay_3114__variable_2417 <= __delay_data_3114__variable_2417;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3118__delay_3117_reinterpretcast_2432 <= __delay_data_3117_reinterpretcast_2432;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _cond_data_2434 <= (_pointer_data_2424)? -17'sd32768 : __delay_data_3110__delay_3109_reinterpretcast_2428;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _cond_data_2439 <= (_pointer_data_2424)? -17'sd32768 : __delay_data_3118__delay_3117_reinterpretcast_2432;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3113__delay_3112__delay_3111__variable_2420 <= __delay_data_3112__delay_3111__variable_2420;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_3116__delay_3115__delay_3114__variable_2417 <= __delay_data_3115__delay_3114__variable_2417;
      end 
      if(_set_flag_2053) begin
        _stream_max_pool_serial_6_parameter_0_next_parameter_data <= 4;
      end 
      if(_stream_max_pool_serial_6_source_start) begin
        __variable_wdata_2417 <= _stream_max_pool_serial_6_parameter_0_next_parameter_data;
      end 
      if(_set_flag_2054) begin
        _stream_max_pool_serial_6_parameter_2_next_parameter_data <= max_pool_serial_6_stream_pad_masks;
      end 
      if(_stream_max_pool_serial_6_source_start) begin
        __variable_wdata_2419 <= _stream_max_pool_serial_6_parameter_2_next_parameter_data;
      end 
      if(_set_flag_2055) begin
        _stream_max_pool_serial_6_source_1_source_mode <= 5'b10;
        _stream_max_pool_serial_6_source_1_source_offset <= max_pool_serial_6_stream_act_local + max_pool_serial_6_act_page_comp_offset_buf;
      end 
      if(_set_flag_2055) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_0 <= 2;
        _source_stream_max_pool_serial_6_source_1_pat_stride_0 <= cparam_max_pool_serial_6_act_read_block;
      end 
      if(_set_flag_2055) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_1 <= 2;
        _source_stream_max_pool_serial_6_source_1_pat_stride_1 <= cparam_max_pool_serial_6_act_read_size;
      end 
      if(_set_flag_2055) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_2 <= cparam_max_pool_serial_6_stream_size;
        _source_stream_max_pool_serial_6_source_1_pat_stride_2 <= 1;
      end 
      if(_set_flag_2055) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_3 <= 1;
        _source_stream_max_pool_serial_6_source_1_pat_stride_3 <= 0;
      end 
      if(_set_flag_2055) begin
        _stream_max_pool_serial_6_source_1_source_sel <= 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_offset_buf <= _stream_max_pool_serial_6_source_1_source_offset;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_0 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_1 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_2 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_3 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_2;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_3;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0 <= _source_stream_max_pool_serial_6_source_1_pat_stride_0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1 <= _source_stream_max_pool_serial_6_source_1_pat_stride_1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2 <= _source_stream_max_pool_serial_6_source_1_pat_stride_2;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3 <= _source_stream_max_pool_serial_6_source_1_pat_stride_3;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_busy && _stream_max_pool_serial_6_is_root) begin
        __variable_wdata_2418 <= _stream_max_pool_serial_6_source_1_source_ram_rdata;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_idle <= 0;
        _stream_max_pool_serial_6_source_1_source_ram_raddr <= _stream_max_pool_serial_6_source_1_source_pat_all_offset;
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0;
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_count_0 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1;
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_count_1 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0)) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2;
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_count_2 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0)) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0)) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3;
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_count_3 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0)) && (_source_stream_max_pool_serial_6_source_1_pat_count_3 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_source_stop && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_idle <= 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 2) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_idle <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2059 <= _set_flag_2058;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2060 <= _tmp_2059;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2061 <= _tmp_2060;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2062 <= _tmp_2061;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2063 <= _tmp_2062;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2064 <= _tmp_2063;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2065 <= _tmp_2064;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2068 <= _tmp_2067;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2069 <= _tmp_2068;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2070 <= _tmp_2069;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2071 <= _tmp_2070;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2072 <= _tmp_2071;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2073 <= _tmp_2072;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2074 <= _tmp_2073;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2075 <= cparam_max_pool_serial_6_stream_size;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2076 <= _tmp_2075;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2077 <= _tmp_2076;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2078 <= _tmp_2077;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2079 <= _tmp_2078;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2080 <= _tmp_2079;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2081 <= _tmp_2080;
      end 
      if(_tmp_2065) begin
        _stream_max_pool_serial_6_sink_6_sink_mode <= 5'b1;
        _stream_max_pool_serial_6_sink_6_sink_offset <= _tmp_2074;
        _stream_max_pool_serial_6_sink_6_sink_size <= _tmp_2081;
        _stream_max_pool_serial_6_sink_6_sink_stride <= 1;
      end 
      if(_tmp_2065) begin
        _stream_max_pool_serial_6_sink_6_sink_sel <= 2;
      end 
      if(_stream_max_pool_serial_6_sink_start && _stream_max_pool_serial_6_sink_6_sink_mode & 5'b1 && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_offset_buf <= _stream_max_pool_serial_6_sink_6_sink_offset;
        _stream_max_pool_serial_6_sink_6_sink_size_buf <= _stream_max_pool_serial_6_sink_6_sink_size;
        _stream_max_pool_serial_6_sink_6_sink_stride_buf <= _stream_max_pool_serial_6_sink_6_sink_stride;
      end 
      if((_stream_max_pool_serial_6_sink_6_sink_fsm_1 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_waddr <= _stream_max_pool_serial_6_sink_6_sink_offset_buf - _stream_max_pool_serial_6_sink_6_sink_stride_buf;
        _stream_max_pool_serial_6_sink_6_sink_count <= _stream_max_pool_serial_6_sink_6_sink_size_buf;
      end 
      if((_stream_max_pool_serial_6_sink_6_sink_fsm_1 == 2) && stream_max_pool_serial_6_sink_7_data && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_waddr <= _stream_max_pool_serial_6_sink_6_sink_waddr + _stream_max_pool_serial_6_sink_6_sink_stride_buf;
        _stream_max_pool_serial_6_sink_6_sink_wdata <= stream_max_pool_serial_6_sink_6_data;
        _stream_max_pool_serial_6_sink_6_sink_wenable <= 1;
        _stream_max_pool_serial_6_sink_6_sink_count <= _stream_max_pool_serial_6_sink_6_sink_count - 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2123 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2124 <= _tmp_2123;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2125 <= _tmp_2124;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2126 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2127 <= _tmp_2126;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2128 <= _tmp_2127;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_2128) begin
        __variable_wdata_2420 <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2129 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2130 <= _tmp_2129;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2131 <= _tmp_2130;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2132 <= _tmp_2131;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_2132) begin
        __variable_wdata_2420 <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2135 <= _tmp_2134;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2138 <= _tmp_2137;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_2138) begin
        __variable_wdata_2420 <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2139 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2140 <= _tmp_2139;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2141 <= _tmp_2140;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2142 <= _tmp_2141;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2143 <= _tmp_2142;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2144 <= _tmp_2143;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2145 <= _tmp_2144;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2146 <= _stream_max_pool_serial_6_source_stop;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2147 <= _tmp_2146;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2148 <= _tmp_2147;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2149 <= _tmp_2148;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2150 <= _tmp_2149;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2151 <= _tmp_2150;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2152 <= _tmp_2151;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2153 <= _stream_max_pool_serial_6_source_busy;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2154 <= _tmp_2153;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2155 <= _tmp_2154;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2156 <= _tmp_2155;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2157 <= _tmp_2156;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2158 <= _tmp_2157;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2159 <= _tmp_2158;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_2160 <= _stream_max_pool_serial_6_sink_busy;
      end 
      if(!_stream_max_pool_serial_6_sink_busy && _tmp_2160) begin
        _stream_max_pool_serial_6_busy_reg <= 0;
      end 
      if(_stream_max_pool_serial_6_source_busy) begin
        _stream_max_pool_serial_6_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_max_pool_serial_6_fsm_1 = 1;
  localparam _stream_max_pool_serial_6_fsm_2 = 2;
  localparam _stream_max_pool_serial_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_init;
      _stream_max_pool_serial_6_source_start <= 0;
      _stream_max_pool_serial_6_source_busy <= 0;
      _stream_max_pool_serial_6_stream_ivalid <= 0;
    end else begin
      if(_stream_max_pool_serial_6_stream_oready && _tmp_2125) begin
        _stream_max_pool_serial_6_stream_ivalid <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_2135) begin
        _stream_max_pool_serial_6_stream_ivalid <= 0;
      end 
      case(_stream_max_pool_serial_6_fsm)
        _stream_max_pool_serial_6_fsm_init: begin
          if(_stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_source_start <= 1;
          end 
          if(_stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_1;
          end 
        end
        _stream_max_pool_serial_6_fsm_1: begin
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_start <= 0;
            _stream_max_pool_serial_6_source_busy <= 1;
          end 
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_2;
          end 
        end
        _stream_max_pool_serial_6_fsm_2: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_3;
          end 
        end
        _stream_max_pool_serial_6_fsm_3: begin
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3))) begin
            _stream_max_pool_serial_6_source_busy <= 0;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3)) && _stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_source_start <= 1;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3))) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_init;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3)) && _stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_source_7_source_ram_renable <= 0;
      _stream_matmul_16_source_7_source_fifo_deq <= 0;
      _stream_matmul_16_source_7_idle <= 1;
      _stream_matmul_16_source_9_source_ram_renable <= 0;
      _stream_matmul_16_source_9_source_fifo_deq <= 0;
      _stream_matmul_16_source_9_idle <= 1;
      _stream_matmul_16_source_11_source_ram_renable <= 0;
      _stream_matmul_16_source_11_source_fifo_deq <= 0;
      _stream_matmul_16_source_11_idle <= 1;
      _stream_matmul_16_source_13_source_ram_renable <= 0;
      _stream_matmul_16_source_13_source_fifo_deq <= 0;
      _stream_matmul_16_source_13_idle <= 1;
      _stream_matmul_16_source_15_source_ram_renable <= 0;
      _stream_matmul_16_source_15_source_fifo_deq <= 0;
      _stream_matmul_16_source_15_idle <= 1;
      _stream_matmul_16_source_20_source_ram_renable <= 0;
      _stream_matmul_16_source_20_source_fifo_deq <= 0;
      _stream_matmul_16_source_20_idle <= 1;
      _stream_matmul_16_source_21_source_ram_renable <= 0;
      _stream_matmul_16_source_21_source_fifo_deq <= 0;
      _stream_matmul_16_source_21_idle <= 1;
      _stream_matmul_16_source_22_source_ram_renable <= 0;
      _stream_matmul_16_source_22_source_fifo_deq <= 0;
      _stream_matmul_16_source_22_idle <= 1;
      _stream_matmul_16_sink_33_sink_wenable <= 0;
      _stream_matmul_16_sink_33_sink_fifo_enq <= 0;
      _stream_matmul_16_sink_34_sink_wenable <= 0;
      _stream_matmul_16_sink_34_sink_fifo_enq <= 0;
      __stream_matmul_16_stream_ivalid_1 <= 0;
      __stream_matmul_16_stream_ivalid_2 <= 0;
      __stream_matmul_16_stream_ivalid_3 <= 0;
      __stream_matmul_16_stream_ivalid_4 <= 0;
      __stream_matmul_16_stream_ivalid_5 <= 0;
      __stream_matmul_16_stream_ivalid_6 <= 0;
      __stream_matmul_16_stream_ivalid_7 <= 0;
      __stream_matmul_16_stream_ivalid_8 <= 0;
      __stream_matmul_16_stream_ivalid_9 <= 0;
      __stream_matmul_16_stream_ivalid_10 <= 0;
      __stream_matmul_16_stream_ivalid_11 <= 0;
      __stream_matmul_16_stream_ivalid_12 <= 0;
      __stream_matmul_16_stream_ivalid_13 <= 0;
      __stream_matmul_16_stream_ivalid_14 <= 0;
      __stream_matmul_16_stream_ivalid_15 <= 0;
      __stream_matmul_16_stream_ivalid_16 <= 0;
      __stream_matmul_16_stream_ivalid_17 <= 0;
      __stream_matmul_16_stream_ivalid_18 <= 0;
      __stream_matmul_16_stream_ivalid_19 <= 0;
      __stream_matmul_16_stream_ivalid_20 <= 0;
      __stream_matmul_16_stream_ivalid_21 <= 0;
      __stream_matmul_16_stream_ivalid_22 <= 0;
      __stream_matmul_16_stream_ivalid_23 <= 0;
      __stream_matmul_16_stream_ivalid_24 <= 0;
      __stream_matmul_16_stream_ivalid_25 <= 0;
      __stream_matmul_16_stream_ivalid_26 <= 0;
      __stream_matmul_16_stream_ivalid_27 <= 0;
      __stream_matmul_16_stream_ivalid_28 <= 0;
      __stream_matmul_16_stream_ivalid_29 <= 0;
      __stream_matmul_16_stream_ivalid_30 <= 0;
      __stream_matmul_16_stream_ivalid_31 <= 0;
      __stream_matmul_16_stream_ivalid_32 <= 0;
      _counter_data_2451 <= 1'sd0;
      _counter_count_2451 <= 1'sd0;
      _minus_data_2456 <= 0;
      _minus_data_2462 <= 0;
      _eq_data_2531 <= 0;
      _eq_data_2535 <= 0;
      _plus_data_2582 <= 0;
      _plus_data_2587 <= 0;
      _plus_data_2592 <= 0;
      _plus_data_2597 <= 0;
      _eq_data_2603 <= 0;
      _eq_data_2606 <= 0;
      _plus_data_2613 <= 0;
      _plus_data_2618 <= 0;
      _plus_data_2623 <= 0;
      _plus_data_2628 <= 0;
      _eq_data_2634 <= 0;
      _eq_data_2637 <= 0;
      __delay_data_3119_pointer_2454 <= 0;
      __delay_data_3121__variable_2530 <= 0;
      __delay_data_3124_pointer_2577 <= 0;
      __delay_data_3127_reinterpretcast_2556 <= 0;
      __delay_data_3132_pointer_2460 <= 0;
      __delay_data_3136_reinterpretcast_2560 <= 0;
      __delay_data_3141__variable_2450 <= 0;
      __delay_data_3168__variable_2445 <= 0;
      __delay_data_3182_reinterpretcast_2568 <= 0;
      __delay_data_3187_reinterpretcast_2572 <= 0;
      __delay_data_3205_cond_2477 <= 0;
      __delay_data_3225_cond_2489 <= 0;
      __delay_data_3330_cond_2476 <= 0;
      __delay_data_3350_cond_2488 <= 0;
      _eq_data_2458 <= 0;
      _eq_data_2464 <= 0;
      __delay_data_3120__delay_3119_pointer_2454 <= 0;
      __delay_data_3122_reinterpretcast_2542 <= 0;
      __delay_data_3125__delay_3124_pointer_2577 <= 0;
      __delay_data_3128__delay_3127_reinterpretcast_2556 <= 0;
      __delay_data_3130_plus_2582 <= 0;
      __delay_data_3133__delay_3132_pointer_2460 <= 0;
      __delay_data_3134_reinterpretcast_2546 <= 0;
      __delay_data_3137__delay_3136_reinterpretcast_2560 <= 0;
      __delay_data_3139_plus_2587 <= 0;
      __delay_data_3142__delay_3141__variable_2450 <= 0;
      __delay_data_3155_plus_2592 <= 0;
      __delay_data_3169__delay_3168__variable_2445 <= 0;
      __delay_data_3183__delay_3182_reinterpretcast_2568 <= 0;
      __delay_data_3185_plus_2613 <= 0;
      __delay_data_3188__delay_3187_reinterpretcast_2572 <= 0;
      __delay_data_3190_plus_2618 <= 0;
      __delay_data_3192_plus_2623 <= 0;
      __delay_data_3206__delay_3205_cond_2477 <= 0;
      __delay_data_3226__delay_3225_cond_2489 <= 0;
      __delay_data_3246_plus_2628 <= 0;
      __delay_data_3267_eq_2634 <= 0;
      __delay_data_3299_eq_2637 <= 0;
      __delay_data_3331__delay_3330_cond_2476 <= 0;
      __delay_data_3351__delay_3350_cond_2488 <= 0;
      __delay_data_3371_plus_2597 <= 0;
      __delay_data_3392_eq_2603 <= 0;
      __delay_data_3424_eq_2606 <= 0;
      _land_data_2459 <= 0;
      _land_data_2465 <= 0;
      __delay_data_3123__delay_3122_reinterpretcast_2542 <= 0;
      __delay_data_3126__delay_3125__delay_3124_pointer_2577 <= 0;
      __delay_data_3129__delay_3128__delay_3127_reinterpretcast_2556 <= 0;
      __delay_data_3131__delay_3130_plus_2582 <= 0;
      __delay_data_3135__delay_3134_reinterpretcast_2546 <= 0;
      __delay_data_3138__delay_3137__delay_3136_reinterpretcast_2560 <= 0;
      __delay_data_3140__delay_3139_plus_2587 <= 0;
      __delay_data_3143__delay_3142__delay_3141__variable_2450 <= 0;
      __delay_data_3156__delay_3155_plus_2592 <= 0;
      __delay_data_3170__delay_3169__delay_3168__variable_2445 <= 0;
      __delay_data_3184__delay_3183__delay_3182_reinterpretcast_2568 <= 0;
      __delay_data_3186__delay_3185_plus_2613 <= 0;
      __delay_data_3189__delay_3188__delay_3187_reinterpretcast_2572 <= 0;
      __delay_data_3191__delay_3190_plus_2618 <= 0;
      __delay_data_3193__delay_3192_plus_2623 <= 0;
      __delay_data_3207__delay_3206__delay_3205_cond_2477 <= 0;
      __delay_data_3227__delay_3226__delay_3225_cond_2489 <= 0;
      __delay_data_3247__delay_3246_plus_2628 <= 0;
      __delay_data_3268__delay_3267_eq_2634 <= 0;
      __delay_data_3300__delay_3299_eq_2637 <= 0;
      __delay_data_3332__delay_3331__delay_3330_cond_2476 <= 0;
      __delay_data_3352__delay_3351__delay_3350_cond_2488 <= 0;
      __delay_data_3372__delay_3371_plus_2597 <= 0;
      __delay_data_3393__delay_3392_eq_2603 <= 0;
      __delay_data_3425__delay_3424_eq_2606 <= 0;
      __delay_data_3144__delay_3143__delay_3142____variable_2450 <= 0;
      __delay_data_3157__delay_3156__delay_3155_plus_2592 <= 0;
      __delay_data_3171__delay_3170__delay_3169____variable_2445 <= 0;
      __delay_data_3194__delay_3193__delay_3192_plus_2623 <= 0;
      __delay_data_3208__delay_3207__delay_3206___cond_2477 <= 0;
      __delay_data_3228__delay_3227__delay_3226___cond_2489 <= 0;
      __delay_data_3248__delay_3247__delay_3246_plus_2628 <= 0;
      __delay_data_3269__delay_3268__delay_3267_eq_2634 <= 0;
      __delay_data_3301__delay_3300__delay_3299_eq_2637 <= 0;
      __delay_data_3333__delay_3332__delay_3331___cond_2476 <= 0;
      __delay_data_3353__delay_3352__delay_3351___cond_2488 <= 0;
      __delay_data_3373__delay_3372__delay_3371_plus_2597 <= 0;
      __delay_data_3394__delay_3393__delay_3392_eq_2603 <= 0;
      __delay_data_3426__delay_3425__delay_3424_eq_2606 <= 0;
      __delay_data_3145__delay_3144__delay_3143____variable_2450 <= 0;
      __delay_data_3158__delay_3157__delay_3156___plus_2592 <= 0;
      __delay_data_3172__delay_3171__delay_3170____variable_2445 <= 0;
      __delay_data_3195__delay_3194__delay_3193___plus_2623 <= 0;
      __delay_data_3209__delay_3208__delay_3207___cond_2477 <= 0;
      __delay_data_3229__delay_3228__delay_3227___cond_2489 <= 0;
      __delay_data_3249__delay_3248__delay_3247___plus_2628 <= 0;
      __delay_data_3270__delay_3269__delay_3268__delay_3267_eq_2634 <= 0;
      __delay_data_3302__delay_3301__delay_3300__delay_3299_eq_2637 <= 0;
      __delay_data_3334__delay_3333__delay_3332___cond_2476 <= 0;
      __delay_data_3354__delay_3353__delay_3352___cond_2488 <= 0;
      __delay_data_3374__delay_3373__delay_3372___plus_2597 <= 0;
      __delay_data_3395__delay_3394__delay_3393__delay_3392_eq_2603 <= 0;
      __delay_data_3427__delay_3426__delay_3425__delay_3424_eq_2606 <= 0;
      __delay_data_3146__delay_3145__delay_3144____variable_2450 <= 0;
      __delay_data_3159__delay_3158__delay_3157___plus_2592 <= 0;
      __delay_data_3173__delay_3172__delay_3171____variable_2445 <= 0;
      __delay_data_3196__delay_3195__delay_3194___plus_2623 <= 0;
      __delay_data_3210__delay_3209__delay_3208___cond_2477 <= 0;
      __delay_data_3230__delay_3229__delay_3228___cond_2489 <= 0;
      __delay_data_3250__delay_3249__delay_3248___plus_2628 <= 0;
      __delay_data_3271__delay_3270__delay_3269__delay_3268___eq_2634 <= 0;
      __delay_data_3303__delay_3302__delay_3301__delay_3300___eq_2637 <= 0;
      __delay_data_3335__delay_3334__delay_3333___cond_2476 <= 0;
      __delay_data_3355__delay_3354__delay_3353___cond_2488 <= 0;
      __delay_data_3375__delay_3374__delay_3373___plus_2597 <= 0;
      __delay_data_3396__delay_3395__delay_3394__delay_3393___eq_2603 <= 0;
      __delay_data_3428__delay_3427__delay_3426__delay_3425___eq_2606 <= 0;
      __delay_data_3147__delay_3146__delay_3145____variable_2450 <= 0;
      __delay_data_3160__delay_3159__delay_3158___plus_2592 <= 0;
      __delay_data_3174__delay_3173__delay_3172____variable_2445 <= 0;
      __delay_data_3197__delay_3196__delay_3195___plus_2623 <= 0;
      __delay_data_3211__delay_3210__delay_3209___cond_2477 <= 0;
      __delay_data_3231__delay_3230__delay_3229___cond_2489 <= 0;
      __delay_data_3251__delay_3250__delay_3249___plus_2628 <= 0;
      __delay_data_3272__delay_3271__delay_3270__delay_3269___eq_2634 <= 0;
      __delay_data_3304__delay_3303__delay_3302__delay_3301___eq_2637 <= 0;
      __delay_data_3336__delay_3335__delay_3334___cond_2476 <= 0;
      __delay_data_3356__delay_3355__delay_3354___cond_2488 <= 0;
      __delay_data_3376__delay_3375__delay_3374___plus_2597 <= 0;
      __delay_data_3397__delay_3396__delay_3395__delay_3394___eq_2603 <= 0;
      __delay_data_3429__delay_3428__delay_3427__delay_3426___eq_2606 <= 0;
      __delay_data_3148__delay_3147__delay_3146____variable_2450 <= 0;
      __delay_data_3161__delay_3160__delay_3159___plus_2592 <= 0;
      __delay_data_3175__delay_3174__delay_3173____variable_2445 <= 0;
      __delay_data_3198__delay_3197__delay_3196___plus_2623 <= 0;
      __delay_data_3212__delay_3211__delay_3210___cond_2477 <= 0;
      __delay_data_3232__delay_3231__delay_3230___cond_2489 <= 0;
      __delay_data_3252__delay_3251__delay_3250___plus_2628 <= 0;
      __delay_data_3273__delay_3272__delay_3271__delay_3270___eq_2634 <= 0;
      __delay_data_3305__delay_3304__delay_3303__delay_3302___eq_2637 <= 0;
      __delay_data_3337__delay_3336__delay_3335___cond_2476 <= 0;
      __delay_data_3357__delay_3356__delay_3355___cond_2488 <= 0;
      __delay_data_3377__delay_3376__delay_3375___plus_2597 <= 0;
      __delay_data_3398__delay_3397__delay_3396__delay_3395___eq_2603 <= 0;
      __delay_data_3430__delay_3429__delay_3428__delay_3427___eq_2606 <= 0;
      __delay_data_3149__delay_3148__delay_3147____variable_2450 <= 0;
      __delay_data_3162__delay_3161__delay_3160___plus_2592 <= 0;
      __delay_data_3176__delay_3175__delay_3174____variable_2445 <= 0;
      __delay_data_3199__delay_3198__delay_3197___plus_2623 <= 0;
      __delay_data_3213__delay_3212__delay_3211___cond_2477 <= 0;
      __delay_data_3233__delay_3232__delay_3231___cond_2489 <= 0;
      __delay_data_3253__delay_3252__delay_3251___plus_2628 <= 0;
      __delay_data_3274__delay_3273__delay_3272__delay_3271___eq_2634 <= 0;
      __delay_data_3306__delay_3305__delay_3304__delay_3303___eq_2637 <= 0;
      __delay_data_3338__delay_3337__delay_3336___cond_2476 <= 0;
      __delay_data_3358__delay_3357__delay_3356___cond_2488 <= 0;
      __delay_data_3378__delay_3377__delay_3376___plus_2597 <= 0;
      __delay_data_3399__delay_3398__delay_3397__delay_3396___eq_2603 <= 0;
      __delay_data_3431__delay_3430__delay_3429__delay_3428___eq_2606 <= 0;
      __delay_data_3150__delay_3149__delay_3148____variable_2450 <= 0;
      __delay_data_3163__delay_3162__delay_3161___plus_2592 <= 0;
      __delay_data_3177__delay_3176__delay_3175____variable_2445 <= 0;
      __delay_data_3200__delay_3199__delay_3198___plus_2623 <= 0;
      __delay_data_3214__delay_3213__delay_3212___cond_2477 <= 0;
      __delay_data_3234__delay_3233__delay_3232___cond_2489 <= 0;
      __delay_data_3254__delay_3253__delay_3252___plus_2628 <= 0;
      __delay_data_3275__delay_3274__delay_3273__delay_3272___eq_2634 <= 0;
      __delay_data_3307__delay_3306__delay_3305__delay_3304___eq_2637 <= 0;
      __delay_data_3339__delay_3338__delay_3337___cond_2476 <= 0;
      __delay_data_3359__delay_3358__delay_3357___cond_2488 <= 0;
      __delay_data_3379__delay_3378__delay_3377___plus_2597 <= 0;
      __delay_data_3400__delay_3399__delay_3398__delay_3397___eq_2603 <= 0;
      __delay_data_3432__delay_3431__delay_3430__delay_3429___eq_2606 <= 0;
      __delay_data_3151__delay_3150__delay_3149____variable_2450 <= 0;
      __delay_data_3164__delay_3163__delay_3162___plus_2592 <= 0;
      __delay_data_3178__delay_3177__delay_3176____variable_2445 <= 0;
      __delay_data_3201__delay_3200__delay_3199___plus_2623 <= 0;
      __delay_data_3215__delay_3214__delay_3213___cond_2477 <= 0;
      __delay_data_3235__delay_3234__delay_3233___cond_2489 <= 0;
      __delay_data_3255__delay_3254__delay_3253___plus_2628 <= 0;
      __delay_data_3276__delay_3275__delay_3274__delay_3273___eq_2634 <= 0;
      __delay_data_3308__delay_3307__delay_3306__delay_3305___eq_2637 <= 0;
      __delay_data_3340__delay_3339__delay_3338___cond_2476 <= 0;
      __delay_data_3360__delay_3359__delay_3358___cond_2488 <= 0;
      __delay_data_3380__delay_3379__delay_3378___plus_2597 <= 0;
      __delay_data_3401__delay_3400__delay_3399__delay_3398___eq_2603 <= 0;
      __delay_data_3433__delay_3432__delay_3431__delay_3430___eq_2606 <= 0;
      __delay_data_3152__delay_3151__delay_3150____variable_2450 <= 0;
      __delay_data_3165__delay_3164__delay_3163___plus_2592 <= 0;
      __delay_data_3179__delay_3178__delay_3177____variable_2445 <= 0;
      __delay_data_3202__delay_3201__delay_3200___plus_2623 <= 0;
      __delay_data_3216__delay_3215__delay_3214___cond_2477 <= 0;
      __delay_data_3236__delay_3235__delay_3234___cond_2489 <= 0;
      __delay_data_3256__delay_3255__delay_3254___plus_2628 <= 0;
      __delay_data_3277__delay_3276__delay_3275__delay_3274___eq_2634 <= 0;
      __delay_data_3309__delay_3308__delay_3307__delay_3306___eq_2637 <= 0;
      __delay_data_3341__delay_3340__delay_3339___cond_2476 <= 0;
      __delay_data_3361__delay_3360__delay_3359___cond_2488 <= 0;
      __delay_data_3381__delay_3380__delay_3379___plus_2597 <= 0;
      __delay_data_3402__delay_3401__delay_3400__delay_3399___eq_2603 <= 0;
      __delay_data_3434__delay_3433__delay_3432__delay_3431___eq_2606 <= 0;
      __delay_data_3153__delay_3152__delay_3151____variable_2450 <= 0;
      __delay_data_3166__delay_3165__delay_3164___plus_2592 <= 0;
      __delay_data_3180__delay_3179__delay_3178____variable_2445 <= 0;
      __delay_data_3203__delay_3202__delay_3201___plus_2623 <= 0;
      __delay_data_3217__delay_3216__delay_3215___cond_2477 <= 0;
      __delay_data_3237__delay_3236__delay_3235___cond_2489 <= 0;
      __delay_data_3257__delay_3256__delay_3255___plus_2628 <= 0;
      __delay_data_3278__delay_3277__delay_3276__delay_3275___eq_2634 <= 0;
      __delay_data_3310__delay_3309__delay_3308__delay_3307___eq_2637 <= 0;
      __delay_data_3342__delay_3341__delay_3340___cond_2476 <= 0;
      __delay_data_3362__delay_3361__delay_3360___cond_2488 <= 0;
      __delay_data_3382__delay_3381__delay_3380___plus_2597 <= 0;
      __delay_data_3403__delay_3402__delay_3401__delay_3400___eq_2603 <= 0;
      __delay_data_3435__delay_3434__delay_3433__delay_3432___eq_2606 <= 0;
      __delay_data_3154__delay_3153__delay_3152____variable_2450 <= 0;
      __delay_data_3167__delay_3166__delay_3165___plus_2592 <= 0;
      __delay_data_3181__delay_3180__delay_3179____variable_2445 <= 0;
      __delay_data_3204__delay_3203__delay_3202___plus_2623 <= 0;
      __delay_data_3218__delay_3217__delay_3216___cond_2477 <= 0;
      __delay_data_3238__delay_3237__delay_3236___cond_2489 <= 0;
      __delay_data_3258__delay_3257__delay_3256___plus_2628 <= 0;
      __delay_data_3279__delay_3278__delay_3277__delay_3276___eq_2634 <= 0;
      __delay_data_3311__delay_3310__delay_3309__delay_3308___eq_2637 <= 0;
      __delay_data_3343__delay_3342__delay_3341___cond_2476 <= 0;
      __delay_data_3363__delay_3362__delay_3361___cond_2488 <= 0;
      __delay_data_3383__delay_3382__delay_3381___plus_2597 <= 0;
      __delay_data_3404__delay_3403__delay_3402__delay_3401___eq_2603 <= 0;
      __delay_data_3436__delay_3435__delay_3434__delay_3433___eq_2606 <= 0;
      __delay_data_3219__delay_3218__delay_3217___cond_2477 <= 0;
      __delay_data_3239__delay_3238__delay_3237___cond_2489 <= 0;
      __delay_data_3259__delay_3258__delay_3257___plus_2628 <= 0;
      __delay_data_3280__delay_3279__delay_3278__delay_3277___eq_2634 <= 0;
      __delay_data_3312__delay_3311__delay_3310__delay_3309___eq_2637 <= 0;
      __delay_data_3344__delay_3343__delay_3342___cond_2476 <= 0;
      __delay_data_3364__delay_3363__delay_3362___cond_2488 <= 0;
      __delay_data_3384__delay_3383__delay_3382___plus_2597 <= 0;
      __delay_data_3405__delay_3404__delay_3403__delay_3402___eq_2603 <= 0;
      __delay_data_3437__delay_3436__delay_3435__delay_3434___eq_2606 <= 0;
      __delay_data_3220__delay_3219__delay_3218___cond_2477 <= 0;
      __delay_data_3240__delay_3239__delay_3238___cond_2489 <= 0;
      __delay_data_3260__delay_3259__delay_3258___plus_2628 <= 0;
      __delay_data_3281__delay_3280__delay_3279__delay_3278___eq_2634 <= 0;
      __delay_data_3313__delay_3312__delay_3311__delay_3310___eq_2637 <= 0;
      __delay_data_3345__delay_3344__delay_3343___cond_2476 <= 0;
      __delay_data_3365__delay_3364__delay_3363___cond_2488 <= 0;
      __delay_data_3385__delay_3384__delay_3383___plus_2597 <= 0;
      __delay_data_3406__delay_3405__delay_3404__delay_3403___eq_2603 <= 0;
      __delay_data_3438__delay_3437__delay_3436__delay_3435___eq_2606 <= 0;
      __delay_data_3221__delay_3220__delay_3219___cond_2477 <= 0;
      __delay_data_3241__delay_3240__delay_3239___cond_2489 <= 0;
      __delay_data_3261__delay_3260__delay_3259___plus_2628 <= 0;
      __delay_data_3282__delay_3281__delay_3280__delay_3279___eq_2634 <= 0;
      __delay_data_3314__delay_3313__delay_3312__delay_3311___eq_2637 <= 0;
      __delay_data_3346__delay_3345__delay_3344___cond_2476 <= 0;
      __delay_data_3366__delay_3365__delay_3364___cond_2488 <= 0;
      __delay_data_3386__delay_3385__delay_3384___plus_2597 <= 0;
      __delay_data_3407__delay_3406__delay_3405__delay_3404___eq_2603 <= 0;
      __delay_data_3439__delay_3438__delay_3437__delay_3436___eq_2606 <= 0;
      __delay_data_3222__delay_3221__delay_3220___cond_2477 <= 0;
      __delay_data_3242__delay_3241__delay_3240___cond_2489 <= 0;
      __delay_data_3262__delay_3261__delay_3260___plus_2628 <= 0;
      __delay_data_3283__delay_3282__delay_3281__delay_3280___eq_2634 <= 0;
      __delay_data_3315__delay_3314__delay_3313__delay_3312___eq_2637 <= 0;
      __delay_data_3347__delay_3346__delay_3345___cond_2476 <= 0;
      __delay_data_3367__delay_3366__delay_3365___cond_2488 <= 0;
      __delay_data_3387__delay_3386__delay_3385___plus_2597 <= 0;
      __delay_data_3408__delay_3407__delay_3406__delay_3405___eq_2603 <= 0;
      __delay_data_3440__delay_3439__delay_3438__delay_3437___eq_2606 <= 0;
      __delay_data_3223__delay_3222__delay_3221___cond_2477 <= 0;
      __delay_data_3243__delay_3242__delay_3241___cond_2489 <= 0;
      __delay_data_3263__delay_3262__delay_3261___plus_2628 <= 0;
      __delay_data_3284__delay_3283__delay_3282__delay_3281___eq_2634 <= 0;
      __delay_data_3316__delay_3315__delay_3314__delay_3313___eq_2637 <= 0;
      __delay_data_3348__delay_3347__delay_3346___cond_2476 <= 0;
      __delay_data_3368__delay_3367__delay_3366___cond_2488 <= 0;
      __delay_data_3388__delay_3387__delay_3386___plus_2597 <= 0;
      __delay_data_3409__delay_3408__delay_3407__delay_3406___eq_2603 <= 0;
      __delay_data_3441__delay_3440__delay_3439__delay_3438___eq_2606 <= 0;
      __delay_data_3224__delay_3223__delay_3222___cond_2477 <= 0;
      __delay_data_3244__delay_3243__delay_3242___cond_2489 <= 0;
      __delay_data_3264__delay_3263__delay_3262___plus_2628 <= 0;
      __delay_data_3285__delay_3284__delay_3283__delay_3282___eq_2634 <= 0;
      __delay_data_3317__delay_3316__delay_3315__delay_3314___eq_2637 <= 0;
      __delay_data_3349__delay_3348__delay_3347___cond_2476 <= 0;
      __delay_data_3369__delay_3368__delay_3367___cond_2488 <= 0;
      __delay_data_3389__delay_3388__delay_3387___plus_2597 <= 0;
      __delay_data_3410__delay_3409__delay_3408__delay_3407___eq_2603 <= 0;
      __delay_data_3442__delay_3441__delay_3440__delay_3439___eq_2606 <= 0;
      _plus_data_2595 <= 0;
      _plus_data_2626 <= 0;
      __delay_data_3245__delay_3244__delay_3243___cond_2489 <= 0;
      __delay_data_3265__delay_3264__delay_3263___plus_2628 <= 0;
      __delay_data_3286__delay_3285__delay_3284__delay_3283___eq_2634 <= 0;
      __delay_data_3318__delay_3317__delay_3316__delay_3315___eq_2637 <= 0;
      __delay_data_3370__delay_3369__delay_3368___cond_2488 <= 0;
      __delay_data_3390__delay_3389__delay_3388___plus_2597 <= 0;
      __delay_data_3411__delay_3410__delay_3409__delay_3408___eq_2603 <= 0;
      __delay_data_3443__delay_3442__delay_3441__delay_3440___eq_2606 <= 0;
      __delay_data_3455__substreamoutput_2594 <= 0;
      __delay_data_3287__delay_3286__delay_3285__delay_3284___eq_2634 <= 0;
      __delay_data_3319__delay_3318__delay_3317__delay_3316___eq_2637 <= 0;
      __delay_data_3412__delay_3411__delay_3410__delay_3409___eq_2603 <= 0;
      __delay_data_3444__delay_3443__delay_3442__delay_3441___eq_2606 <= 0;
      __delay_data_3456__delay_3455__substreamoutput_2594 <= 0;
      __delay_data_3288__delay_3287__delay_3286__delay_3285___eq_2634 <= 0;
      __delay_data_3320__delay_3319__delay_3318__delay_3317___eq_2637 <= 0;
      __delay_data_3413__delay_3412__delay_3411__delay_3410___eq_2603 <= 0;
      __delay_data_3445__delay_3444__delay_3443__delay_3442___eq_2606 <= 0;
      __delay_data_3457__delay_3456____substreamoutput_2594 <= 0;
      __delay_data_3289__delay_3288__delay_3287__delay_3286___eq_2634 <= 0;
      __delay_data_3321__delay_3320__delay_3319__delay_3318___eq_2637 <= 0;
      __delay_data_3414__delay_3413__delay_3412__delay_3411___eq_2603 <= 0;
      __delay_data_3446__delay_3445__delay_3444__delay_3443___eq_2606 <= 0;
      __delay_data_3458__delay_3457____substreamoutput_2594 <= 0;
      __delay_data_3290__delay_3289__delay_3288__delay_3287___eq_2634 <= 0;
      __delay_data_3322__delay_3321__delay_3320__delay_3319___eq_2637 <= 0;
      __delay_data_3415__delay_3414__delay_3413__delay_3412___eq_2603 <= 0;
      __delay_data_3447__delay_3446__delay_3445__delay_3444___eq_2606 <= 0;
      __delay_data_3459__delay_3458____substreamoutput_2594 <= 0;
      __delay_data_3291__delay_3290__delay_3289__delay_3288___eq_2634 <= 0;
      __delay_data_3323__delay_3322__delay_3321__delay_3320___eq_2637 <= 0;
      __delay_data_3416__delay_3415__delay_3414__delay_3413___eq_2603 <= 0;
      __delay_data_3448__delay_3447__delay_3446__delay_3445___eq_2606 <= 0;
      __delay_data_3460__delay_3459____substreamoutput_2594 <= 0;
      __delay_data_3292__delay_3291__delay_3290__delay_3289___eq_2634 <= 0;
      __delay_data_3324__delay_3323__delay_3322__delay_3321___eq_2637 <= 0;
      __delay_data_3417__delay_3416__delay_3415__delay_3414___eq_2603 <= 0;
      __delay_data_3449__delay_3448__delay_3447__delay_3446___eq_2606 <= 0;
      __delay_data_3461__delay_3460____substreamoutput_2594 <= 0;
      __delay_data_3293__delay_3292__delay_3291__delay_3290___eq_2634 <= 0;
      __delay_data_3325__delay_3324__delay_3323__delay_3322___eq_2637 <= 0;
      __delay_data_3418__delay_3417__delay_3416__delay_3415___eq_2603 <= 0;
      __delay_data_3450__delay_3449__delay_3448__delay_3447___eq_2606 <= 0;
      __delay_data_3462__delay_3461____substreamoutput_2594 <= 0;
      __delay_data_3294__delay_3293__delay_3292__delay_3291___eq_2634 <= 0;
      __delay_data_3326__delay_3325__delay_3324__delay_3323___eq_2637 <= 0;
      __delay_data_3419__delay_3418__delay_3417__delay_3416___eq_2603 <= 0;
      __delay_data_3451__delay_3450__delay_3449__delay_3448___eq_2606 <= 0;
      __delay_data_3463__delay_3462____substreamoutput_2594 <= 0;
      __delay_data_3295__delay_3294__delay_3293__delay_3292___eq_2634 <= 0;
      __delay_data_3327__delay_3326__delay_3325__delay_3324___eq_2637 <= 0;
      __delay_data_3420__delay_3419__delay_3418__delay_3417___eq_2603 <= 0;
      __delay_data_3452__delay_3451__delay_3450__delay_3449___eq_2606 <= 0;
      __delay_data_3464__delay_3463____substreamoutput_2594 <= 0;
      _greaterthan_data_2600 <= 0;
      _greaterthan_data_2631 <= 0;
      __delay_data_3266__substreamoutput_2629 <= 0;
      __delay_data_3296__delay_3295__delay_3294__delay_3293___eq_2634 <= 0;
      __delay_data_3328__delay_3327__delay_3326__delay_3325___eq_2637 <= 0;
      __delay_data_3391__substreamoutput_2598 <= 0;
      __delay_data_3421__delay_3420__delay_3419__delay_3418___eq_2603 <= 0;
      __delay_data_3453__delay_3452__delay_3451__delay_3450___eq_2606 <= 0;
      __delay_data_3465__delay_3464____substreamoutput_2594 <= 0;
      _cond_data_2602 <= 0;
      _cond_data_2633 <= 0;
      __delay_data_3297__delay_3296__delay_3295__delay_3294___eq_2634 <= 0;
      __delay_data_3298__delay_3266__substreamoutput_2629 <= 0;
      __delay_data_3329__delay_3328__delay_3327__delay_3326___eq_2637 <= 0;
      __delay_data_3422__delay_3421__delay_3420__delay_3419___eq_2603 <= 0;
      __delay_data_3423__delay_3391__substreamoutput_2598 <= 0;
      __delay_data_3454__delay_3453__delay_3452__delay_3451___eq_2606 <= 0;
      __delay_data_3466__delay_3465____substreamoutput_2594 <= 0;
      _stream_matmul_16_parameter_0_next_parameter_data <= 0;
      __variable_wdata_2445 <= 0;
      _stream_matmul_16_parameter_1_next_parameter_data <= 0;
      __variable_wdata_2446 <= 0;
      _stream_matmul_16_parameter_2_next_parameter_data <= 0;
      __variable_wdata_2447 <= 0;
      _stream_matmul_16_parameter_3_next_parameter_data <= 0;
      __variable_wdata_2448 <= 0;
      _stream_matmul_16_parameter_4_next_parameter_data <= 0;
      __variable_wdata_2449 <= 0;
      _stream_matmul_16_parameter_6_next_parameter_data <= 0;
      __variable_wdata_2466 <= 0;
      _stream_matmul_16_source_7_source_mode <= 5'b0;
      _stream_matmul_16_source_7_source_offset <= 0;
      _source_stream_matmul_16_source_7_pat_size_0 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_0 <= 0;
      _source_stream_matmul_16_source_7_pat_size_1 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_1 <= 0;
      _source_stream_matmul_16_source_7_pat_size_2 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_2 <= 0;
      _source_stream_matmul_16_source_7_pat_size_3 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_3 <= 0;
      _stream_matmul_16_source_7_source_sel <= 0;
      _stream_matmul_16_source_7_source_offset_buf <= 0;
      _source_stream_matmul_16_source_7_pat_cur_offset_0 <= 0;
      _source_stream_matmul_16_source_7_pat_cur_offset_1 <= 0;
      _source_stream_matmul_16_source_7_pat_cur_offset_2 <= 0;
      _source_stream_matmul_16_source_7_pat_cur_offset_3 <= 0;
      _source_stream_matmul_16_source_7_pat_count_0 <= 0;
      _source_stream_matmul_16_source_7_pat_count_1 <= 0;
      _source_stream_matmul_16_source_7_pat_count_2 <= 0;
      _source_stream_matmul_16_source_7_pat_count_3 <= 0;
      _source_stream_matmul_16_source_7_pat_size_buf_0 <= 0;
      _source_stream_matmul_16_source_7_pat_size_buf_1 <= 0;
      _source_stream_matmul_16_source_7_pat_size_buf_2 <= 0;
      _source_stream_matmul_16_source_7_pat_size_buf_3 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_buf_0 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_buf_1 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_buf_2 <= 0;
      _source_stream_matmul_16_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_2467 <= 0;
      _stream_matmul_16_source_7_source_ram_raddr <= 0;
      _stream_matmul_16_parameter_8_next_parameter_data <= 0;
      __variable_wdata_2478 <= 0;
      _stream_matmul_16_source_9_source_mode <= 5'b0;
      _stream_matmul_16_source_9_source_offset <= 0;
      _source_stream_matmul_16_source_9_pat_size_0 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_0 <= 0;
      _source_stream_matmul_16_source_9_pat_size_1 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_1 <= 0;
      _source_stream_matmul_16_source_9_pat_size_2 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_2 <= 0;
      _source_stream_matmul_16_source_9_pat_size_3 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_3 <= 0;
      _stream_matmul_16_source_9_source_sel <= 0;
      _stream_matmul_16_source_9_source_offset_buf <= 0;
      _source_stream_matmul_16_source_9_pat_cur_offset_0 <= 0;
      _source_stream_matmul_16_source_9_pat_cur_offset_1 <= 0;
      _source_stream_matmul_16_source_9_pat_cur_offset_2 <= 0;
      _source_stream_matmul_16_source_9_pat_cur_offset_3 <= 0;
      _source_stream_matmul_16_source_9_pat_count_0 <= 0;
      _source_stream_matmul_16_source_9_pat_count_1 <= 0;
      _source_stream_matmul_16_source_9_pat_count_2 <= 0;
      _source_stream_matmul_16_source_9_pat_count_3 <= 0;
      _source_stream_matmul_16_source_9_pat_size_buf_0 <= 0;
      _source_stream_matmul_16_source_9_pat_size_buf_1 <= 0;
      _source_stream_matmul_16_source_9_pat_size_buf_2 <= 0;
      _source_stream_matmul_16_source_9_pat_size_buf_3 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_buf_0 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_buf_1 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_buf_2 <= 0;
      _source_stream_matmul_16_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_2479 <= 0;
      _stream_matmul_16_source_9_source_ram_raddr <= 0;
      _stream_matmul_16_parameter_10_next_parameter_data <= 0;
      __variable_wdata_2490 <= 0;
      _stream_matmul_16_source_11_source_mode <= 5'b0;
      _stream_matmul_16_source_11_source_empty_data <= 0;
      __variable_wdata_2491 <= 0;
      _stream_matmul_16_parameter_12_next_parameter_data <= 0;
      __variable_wdata_2502 <= 0;
      _stream_matmul_16_source_13_source_mode <= 5'b0;
      _stream_matmul_16_source_13_source_empty_data <= 0;
      __variable_wdata_2503 <= 0;
      _stream_matmul_16_parameter_14_next_parameter_data <= 0;
      __variable_wdata_2514 <= 0;
      _stream_matmul_16_source_15_source_mode <= 5'b0;
      _stream_matmul_16_source_15_source_empty_data <= 0;
      __variable_wdata_2515 <= 0;
      _stream_matmul_16_parameter_16_next_parameter_data <= 0;
      __variable_wdata_2526 <= 0;
      _stream_matmul_16_parameter_17_next_parameter_data <= 0;
      __variable_wdata_2527 <= 0;
      _stream_matmul_16_parameter_18_next_parameter_data <= 0;
      __variable_wdata_2528 <= 0;
      _stream_matmul_16_parameter_19_next_parameter_data <= 0;
      __variable_wdata_2529 <= 0;
      _stream_matmul_16_source_20_source_mode <= 5'b0;
      _stream_matmul_16_source_20_source_offset <= 0;
      _source_stream_matmul_16_source_20_pat_size_0 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_0 <= 0;
      _source_stream_matmul_16_source_20_pat_size_1 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_1 <= 0;
      _source_stream_matmul_16_source_20_pat_size_2 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_2 <= 0;
      _source_stream_matmul_16_source_20_pat_size_3 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_3 <= 0;
      _stream_matmul_16_source_20_source_sel <= 0;
      _stream_matmul_16_source_20_source_offset_buf <= 0;
      _source_stream_matmul_16_source_20_pat_cur_offset_0 <= 0;
      _source_stream_matmul_16_source_20_pat_cur_offset_1 <= 0;
      _source_stream_matmul_16_source_20_pat_cur_offset_2 <= 0;
      _source_stream_matmul_16_source_20_pat_cur_offset_3 <= 0;
      _source_stream_matmul_16_source_20_pat_count_0 <= 0;
      _source_stream_matmul_16_source_20_pat_count_1 <= 0;
      _source_stream_matmul_16_source_20_pat_count_2 <= 0;
      _source_stream_matmul_16_source_20_pat_count_3 <= 0;
      _source_stream_matmul_16_source_20_pat_size_buf_0 <= 0;
      _source_stream_matmul_16_source_20_pat_size_buf_1 <= 0;
      _source_stream_matmul_16_source_20_pat_size_buf_2 <= 0;
      _source_stream_matmul_16_source_20_pat_size_buf_3 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_buf_0 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_buf_1 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_buf_2 <= 0;
      _source_stream_matmul_16_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_2530 <= 0;
      _stream_matmul_16_source_20_source_ram_raddr <= 0;
      _stream_matmul_16_source_21_source_mode <= 5'b0;
      _stream_matmul_16_source_21_source_offset <= 0;
      _source_stream_matmul_16_source_21_pat_size_0 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_0 <= 0;
      _source_stream_matmul_16_source_21_pat_size_1 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_1 <= 0;
      _source_stream_matmul_16_source_21_pat_size_2 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_2 <= 0;
      _source_stream_matmul_16_source_21_pat_size_3 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_3 <= 0;
      _stream_matmul_16_source_21_source_sel <= 0;
      _stream_matmul_16_source_21_source_offset_buf <= 0;
      _source_stream_matmul_16_source_21_pat_cur_offset_0 <= 0;
      _source_stream_matmul_16_source_21_pat_cur_offset_1 <= 0;
      _source_stream_matmul_16_source_21_pat_cur_offset_2 <= 0;
      _source_stream_matmul_16_source_21_pat_cur_offset_3 <= 0;
      _source_stream_matmul_16_source_21_pat_count_0 <= 0;
      _source_stream_matmul_16_source_21_pat_count_1 <= 0;
      _source_stream_matmul_16_source_21_pat_count_2 <= 0;
      _source_stream_matmul_16_source_21_pat_count_3 <= 0;
      _source_stream_matmul_16_source_21_pat_size_buf_0 <= 0;
      _source_stream_matmul_16_source_21_pat_size_buf_1 <= 0;
      _source_stream_matmul_16_source_21_pat_size_buf_2 <= 0;
      _source_stream_matmul_16_source_21_pat_size_buf_3 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_buf_0 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_buf_1 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_buf_2 <= 0;
      _source_stream_matmul_16_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_2551 <= 0;
      _stream_matmul_16_source_21_source_ram_raddr <= 0;
      _stream_matmul_16_source_22_source_mode <= 5'b0;
      _stream_matmul_16_source_22_source_offset <= 0;
      _source_stream_matmul_16_source_22_pat_size_0 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_0 <= 0;
      _source_stream_matmul_16_source_22_pat_size_1 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_1 <= 0;
      _source_stream_matmul_16_source_22_pat_size_2 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_2 <= 0;
      _source_stream_matmul_16_source_22_pat_size_3 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_3 <= 0;
      _stream_matmul_16_source_22_source_sel <= 0;
      _stream_matmul_16_source_22_source_offset_buf <= 0;
      _source_stream_matmul_16_source_22_pat_cur_offset_0 <= 0;
      _source_stream_matmul_16_source_22_pat_cur_offset_1 <= 0;
      _source_stream_matmul_16_source_22_pat_cur_offset_2 <= 0;
      _source_stream_matmul_16_source_22_pat_cur_offset_3 <= 0;
      _source_stream_matmul_16_source_22_pat_count_0 <= 0;
      _source_stream_matmul_16_source_22_pat_count_1 <= 0;
      _source_stream_matmul_16_source_22_pat_count_2 <= 0;
      _source_stream_matmul_16_source_22_pat_count_3 <= 0;
      _source_stream_matmul_16_source_22_pat_size_buf_0 <= 0;
      _source_stream_matmul_16_source_22_pat_size_buf_1 <= 0;
      _source_stream_matmul_16_source_22_pat_size_buf_2 <= 0;
      _source_stream_matmul_16_source_22_pat_size_buf_3 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_buf_0 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_buf_1 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_buf_2 <= 0;
      _source_stream_matmul_16_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_2552 <= 0;
      _stream_matmul_16_source_22_source_ram_raddr <= 0;
      _tmp_2240 <= 0;
      _tmp_2241 <= 0;
      _tmp_2242 <= 0;
      _tmp_2243 <= 0;
      _tmp_2244 <= 0;
      _tmp_2245 <= 0;
      _tmp_2246 <= 0;
      _tmp_2247 <= 0;
      _tmp_2248 <= 0;
      _tmp_2249 <= 0;
      _tmp_2250 <= 0;
      _tmp_2251 <= 0;
      _tmp_2252 <= 0;
      _tmp_2253 <= 0;
      _tmp_2254 <= 0;
      _tmp_2255 <= 0;
      _tmp_2256 <= 0;
      _tmp_2257 <= 0;
      _tmp_2258 <= 0;
      _tmp_2259 <= 0;
      _tmp_2260 <= 0;
      _tmp_2261 <= 0;
      _tmp_2262 <= 0;
      _tmp_2263 <= 0;
      _tmp_2264 <= 0;
      _tmp_2265 <= 0;
      _tmp_2266 <= 0;
      _tmp_2267 <= 0;
      _tmp_2268 <= 0;
      _tmp_2269 <= 0;
      _tmp_2270 <= 0;
      _tmp_2271 <= 0;
      _tmp_2272 <= 0;
      _tmp_2273 <= 0;
      _tmp_2276 <= 0;
      _tmp_2277 <= 0;
      _tmp_2278 <= 0;
      _tmp_2279 <= 0;
      _tmp_2280 <= 0;
      _tmp_2281 <= 0;
      _tmp_2282 <= 0;
      _tmp_2283 <= 0;
      _tmp_2284 <= 0;
      _tmp_2285 <= 0;
      _tmp_2286 <= 0;
      _tmp_2287 <= 0;
      _tmp_2288 <= 0;
      _tmp_2289 <= 0;
      _tmp_2290 <= 0;
      _tmp_2291 <= 0;
      _tmp_2292 <= 0;
      _tmp_2293 <= 0;
      _tmp_2294 <= 0;
      _tmp_2295 <= 0;
      _tmp_2296 <= 0;
      _tmp_2297 <= 0;
      _tmp_2298 <= 0;
      _tmp_2299 <= 0;
      _tmp_2300 <= 0;
      _tmp_2301 <= 0;
      _tmp_2302 <= 0;
      _tmp_2303 <= 0;
      _tmp_2304 <= 0;
      _tmp_2305 <= 0;
      _tmp_2306 <= 0;
      _tmp_2307 <= 0;
      _tmp_2308 <= 0;
      _tmp_2309 <= 0;
      _tmp_2310 <= 0;
      _tmp_2311 <= 0;
      _tmp_2312 <= 0;
      _tmp_2313 <= 0;
      _tmp_2314 <= 0;
      _tmp_2315 <= 0;
      _tmp_2316 <= 0;
      _tmp_2317 <= 0;
      _tmp_2318 <= 0;
      _tmp_2319 <= 0;
      _tmp_2320 <= 0;
      _tmp_2321 <= 0;
      _tmp_2322 <= 0;
      _tmp_2323 <= 0;
      _tmp_2324 <= 0;
      _tmp_2325 <= 0;
      _tmp_2326 <= 0;
      _tmp_2327 <= 0;
      _tmp_2328 <= 0;
      _tmp_2329 <= 0;
      _tmp_2330 <= 0;
      _tmp_2331 <= 0;
      _tmp_2332 <= 0;
      _tmp_2333 <= 0;
      _tmp_2334 <= 0;
      _tmp_2335 <= 0;
      _tmp_2336 <= 0;
      _tmp_2337 <= 0;
      _tmp_2338 <= 0;
      _tmp_2339 <= 0;
      _tmp_2340 <= 0;
      _tmp_2341 <= 0;
      _tmp_2342 <= 0;
      _tmp_2343 <= 0;
      _stream_matmul_16_sink_33_sink_mode <= 5'b0;
      _stream_matmul_16_sink_33_sink_offset <= 0;
      _stream_matmul_16_sink_33_sink_size <= 0;
      _stream_matmul_16_sink_33_sink_stride <= 0;
      _stream_matmul_16_sink_33_sink_sel <= 0;
      _stream_matmul_16_sink_33_sink_offset_buf <= 0;
      _stream_matmul_16_sink_33_sink_size_buf <= 0;
      _stream_matmul_16_sink_33_sink_stride_buf <= 0;
      _stream_matmul_16_sink_33_sink_waddr <= 0;
      _stream_matmul_16_sink_33_sink_count <= 0;
      _stream_matmul_16_sink_33_sink_wdata <= 0;
      _tmp_2371 <= 0;
      _tmp_2372 <= 0;
      _tmp_2373 <= 0;
      _tmp_2374 <= 0;
      _tmp_2375 <= 0;
      _tmp_2376 <= 0;
      __variable_wdata_2450 <= 0;
      _tmp_2377 <= 0;
      _tmp_2378 <= 0;
      _tmp_2379 <= 0;
      _tmp_2380 <= 0;
      _tmp_2383 <= 0;
      _tmp_2386 <= 0;
      _tmp_2387 <= 0;
      _tmp_2388 <= 0;
      _tmp_2389 <= 0;
      _tmp_2390 <= 0;
      _tmp_2391 <= 0;
      _tmp_2392 <= 0;
      _tmp_2393 <= 0;
      _tmp_2394 <= 0;
      _tmp_2395 <= 0;
      _tmp_2396 <= 0;
      _tmp_2397 <= 0;
      _tmp_2398 <= 0;
      _tmp_2399 <= 0;
      _tmp_2400 <= 0;
      _tmp_2401 <= 0;
      _tmp_2402 <= 0;
      _tmp_2403 <= 0;
      _tmp_2404 <= 0;
      _tmp_2405 <= 0;
      _tmp_2406 <= 0;
      _tmp_2407 <= 0;
      _tmp_2408 <= 0;
      _tmp_2409 <= 0;
      _tmp_2410 <= 0;
      _tmp_2411 <= 0;
      _tmp_2412 <= 0;
      _tmp_2413 <= 0;
      _tmp_2414 <= 0;
      _tmp_2415 <= 0;
      _tmp_2416 <= 0;
      _tmp_2417 <= 0;
      _tmp_2418 <= 0;
      _tmp_2419 <= 0;
      _tmp_2420 <= 0;
      _tmp_2421 <= 0;
      _tmp_2422 <= 0;
      _tmp_2423 <= 0;
      _tmp_2424 <= 0;
      _tmp_2425 <= 0;
      _tmp_2426 <= 0;
      _tmp_2427 <= 0;
      _tmp_2428 <= 0;
      _tmp_2429 <= 0;
      _tmp_2430 <= 0;
      _tmp_2431 <= 0;
      _tmp_2432 <= 0;
      _tmp_2433 <= 0;
      _tmp_2434 <= 0;
      _tmp_2435 <= 0;
      _tmp_2436 <= 0;
      _tmp_2437 <= 0;
      _tmp_2438 <= 0;
      _tmp_2439 <= 0;
      _tmp_2440 <= 0;
      _tmp_2441 <= 0;
      _tmp_2442 <= 0;
      _tmp_2443 <= 0;
      _tmp_2444 <= 0;
      _tmp_2445 <= 0;
      _tmp_2446 <= 0;
      _tmp_2447 <= 0;
      _tmp_2448 <= 0;
      _tmp_2449 <= 0;
      _tmp_2450 <= 0;
      _tmp_2451 <= 0;
      _tmp_2452 <= 0;
      _tmp_2453 <= 0;
      _tmp_2454 <= 0;
      _tmp_2455 <= 0;
      _tmp_2456 <= 0;
      _tmp_2457 <= 0;
      _tmp_2458 <= 0;
      _tmp_2459 <= 0;
      _tmp_2460 <= 0;
      _tmp_2461 <= 0;
      _tmp_2462 <= 0;
      _tmp_2463 <= 0;
      _tmp_2464 <= 0;
      _tmp_2465 <= 0;
      _tmp_2466 <= 0;
      _tmp_2467 <= 0;
      _tmp_2468 <= 0;
      _tmp_2469 <= 0;
      _tmp_2470 <= 0;
      _tmp_2471 <= 0;
      _tmp_2472 <= 0;
      _tmp_2473 <= 0;
      _tmp_2474 <= 0;
      _tmp_2475 <= 0;
      _tmp_2476 <= 0;
      _tmp_2477 <= 0;
      _tmp_2478 <= 0;
      _tmp_2479 <= 0;
      _tmp_2480 <= 0;
      _tmp_2481 <= 0;
      _tmp_2482 <= 0;
      _tmp_2483 <= 0;
      _tmp_2484 <= 0;
      _tmp_2485 <= 0;
      _tmp_2486 <= 0;
      _tmp_2487 <= 0;
      _tmp_2488 <= 0;
      _tmp_2489 <= 0;
      _stream_matmul_16_busy_reg <= 0;
    end else begin
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_7_source_ram_renable <= 0;
        _stream_matmul_16_source_7_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_7_idle <= _stream_matmul_16_source_7_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_9_source_ram_renable <= 0;
        _stream_matmul_16_source_9_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_9_idle <= _stream_matmul_16_source_9_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_11_source_ram_renable <= 0;
        _stream_matmul_16_source_11_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_11_idle <= _stream_matmul_16_source_11_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_13_source_ram_renable <= 0;
        _stream_matmul_16_source_13_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_13_idle <= _stream_matmul_16_source_13_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_15_source_ram_renable <= 0;
        _stream_matmul_16_source_15_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_15_idle <= _stream_matmul_16_source_15_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_20_source_ram_renable <= 0;
        _stream_matmul_16_source_20_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_20_idle <= _stream_matmul_16_source_20_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_21_source_ram_renable <= 0;
        _stream_matmul_16_source_21_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_21_idle <= _stream_matmul_16_source_21_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_22_source_ram_renable <= 0;
        _stream_matmul_16_source_22_source_fifo_deq <= 0;
      end 
      _stream_matmul_16_source_22_idle <= _stream_matmul_16_source_22_idle;
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_sink_33_sink_wenable <= 0;
        _stream_matmul_16_sink_33_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _stream_matmul_16_sink_34_sink_wenable <= 0;
        _stream_matmul_16_sink_34_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_1 <= _stream_matmul_16_stream_ivalid;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_2 <= __stream_matmul_16_stream_ivalid_1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_3 <= __stream_matmul_16_stream_ivalid_2;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_4 <= __stream_matmul_16_stream_ivalid_3;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_5 <= __stream_matmul_16_stream_ivalid_4;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_6 <= __stream_matmul_16_stream_ivalid_5;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_7 <= __stream_matmul_16_stream_ivalid_6;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_8 <= __stream_matmul_16_stream_ivalid_7;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_9 <= __stream_matmul_16_stream_ivalid_8;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_10 <= __stream_matmul_16_stream_ivalid_9;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_11 <= __stream_matmul_16_stream_ivalid_10;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_12 <= __stream_matmul_16_stream_ivalid_11;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_13 <= __stream_matmul_16_stream_ivalid_12;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_14 <= __stream_matmul_16_stream_ivalid_13;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_15 <= __stream_matmul_16_stream_ivalid_14;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_16 <= __stream_matmul_16_stream_ivalid_15;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_17 <= __stream_matmul_16_stream_ivalid_16;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_18 <= __stream_matmul_16_stream_ivalid_17;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_19 <= __stream_matmul_16_stream_ivalid_18;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_20 <= __stream_matmul_16_stream_ivalid_19;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_21 <= __stream_matmul_16_stream_ivalid_20;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_22 <= __stream_matmul_16_stream_ivalid_21;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_23 <= __stream_matmul_16_stream_ivalid_22;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_24 <= __stream_matmul_16_stream_ivalid_23;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_25 <= __stream_matmul_16_stream_ivalid_24;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_26 <= __stream_matmul_16_stream_ivalid_25;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_27 <= __stream_matmul_16_stream_ivalid_26;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_28 <= __stream_matmul_16_stream_ivalid_27;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_29 <= __stream_matmul_16_stream_ivalid_28;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_30 <= __stream_matmul_16_stream_ivalid_29;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_31 <= __stream_matmul_16_stream_ivalid_30;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __stream_matmul_16_stream_ivalid_32 <= __stream_matmul_16_stream_ivalid_31;
      end 
      if(_stream_matmul_16_stream_ivalid && _stream_matmul_16_stream_oready && _counter_reset_cond_2451) begin
        _counter_data_2451 <= 1'sd0;
      end 
      if(_stream_matmul_16_stream_ivalid && _stream_matmul_16_stream_oready) begin
        _counter_data_2451 <= _counter_current_count_2451;
      end 
      if(_stream_matmul_16_stream_ivalid && _stream_matmul_16_stream_oready) begin
        _counter_count_2451 <= (_counter_current_count_2451 >= stream_matmul_16_parameter_0_data - 2'sd1)? _counter_current_count_2451 + 2'sd1 - stream_matmul_16_parameter_0_data : _counter_current_count_2451 + 2'sd1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _minus_data_2456 <= stream_matmul_16_parameter_0_data - 2'sd1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _minus_data_2462 <= stream_matmul_16_parameter_0_data - 2'sd1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2531 <= stream_matmul_16_parameter_1_data == 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2535 <= stream_matmul_16_parameter_2_data == 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2582 <= _cond_data_2500 + stream_matmul_16_parameter_16_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2587 <= _cond_data_2500 + stream_matmul_16_parameter_16_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2592 <= _cond_data_2512 + stream_matmul_16_parameter_17_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2597 <= _cond_data_2524 + stream_matmul_16_parameter_18_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2603 <= stream_matmul_16_parameter_19_data == 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2606 <= stream_matmul_16_parameter_19_data == 2'sd1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2613 <= _cond_data_2501 + stream_matmul_16_parameter_16_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2618 <= _cond_data_2501 + stream_matmul_16_parameter_16_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2623 <= _cond_data_2513 + stream_matmul_16_parameter_17_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2628 <= _cond_data_2525 + stream_matmul_16_parameter_18_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2634 <= stream_matmul_16_parameter_19_data == 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2637 <= stream_matmul_16_parameter_19_data == 2'sd1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3119_pointer_2454 <= _pointer_data_2454;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3121__variable_2530 <= stream_matmul_16_source_20_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3124_pointer_2577 <= _pointer_data_2577;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3127_reinterpretcast_2556 <= _reinterpretcast_data_2556;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3132_pointer_2460 <= _pointer_data_2460;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3136_reinterpretcast_2560 <= _reinterpretcast_data_2560;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3141__variable_2450 <= stream_matmul_16__reduce_reset_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3168__variable_2445 <= stream_matmul_16_parameter_0_data;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3182_reinterpretcast_2568 <= _reinterpretcast_data_2568;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3187_reinterpretcast_2572 <= _reinterpretcast_data_2572;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3205_cond_2477 <= _cond_data_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3225_cond_2489 <= _cond_data_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3330_cond_2476 <= _cond_data_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3350_cond_2488 <= _cond_data_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2458 <= _counter_data_2451 == _minus_data_2456;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _eq_data_2464 <= _counter_data_2451 == _minus_data_2462;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3120__delay_3119_pointer_2454 <= __delay_data_3119_pointer_2454;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3122_reinterpretcast_2542 <= _reinterpretcast_data_2542;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3125__delay_3124_pointer_2577 <= __delay_data_3124_pointer_2577;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3128__delay_3127_reinterpretcast_2556 <= __delay_data_3127_reinterpretcast_2556;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3130_plus_2582 <= _plus_data_2582;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3133__delay_3132_pointer_2460 <= __delay_data_3132_pointer_2460;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3134_reinterpretcast_2546 <= _reinterpretcast_data_2546;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3137__delay_3136_reinterpretcast_2560 <= __delay_data_3136_reinterpretcast_2560;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3139_plus_2587 <= _plus_data_2587;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3142__delay_3141__variable_2450 <= __delay_data_3141__variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3155_plus_2592 <= _plus_data_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3169__delay_3168__variable_2445 <= __delay_data_3168__variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3183__delay_3182_reinterpretcast_2568 <= __delay_data_3182_reinterpretcast_2568;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3185_plus_2613 <= _plus_data_2613;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3188__delay_3187_reinterpretcast_2572 <= __delay_data_3187_reinterpretcast_2572;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3190_plus_2618 <= _plus_data_2618;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3192_plus_2623 <= _plus_data_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3206__delay_3205_cond_2477 <= __delay_data_3205_cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3226__delay_3225_cond_2489 <= __delay_data_3225_cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3246_plus_2628 <= _plus_data_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3267_eq_2634 <= _eq_data_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3299_eq_2637 <= _eq_data_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3331__delay_3330_cond_2476 <= __delay_data_3330_cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3351__delay_3350_cond_2488 <= __delay_data_3350_cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3371_plus_2597 <= _plus_data_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3392_eq_2603 <= _eq_data_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3424_eq_2606 <= _eq_data_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _land_data_2459 <= __delay_data_3120__delay_3119_pointer_2454 && _eq_data_2458;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _land_data_2465 <= __delay_data_3133__delay_3132_pointer_2460 && _eq_data_2464;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3123__delay_3122_reinterpretcast_2542 <= __delay_data_3122_reinterpretcast_2542;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3126__delay_3125__delay_3124_pointer_2577 <= __delay_data_3125__delay_3124_pointer_2577;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3129__delay_3128__delay_3127_reinterpretcast_2556 <= __delay_data_3128__delay_3127_reinterpretcast_2556;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3131__delay_3130_plus_2582 <= __delay_data_3130_plus_2582;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3135__delay_3134_reinterpretcast_2546 <= __delay_data_3134_reinterpretcast_2546;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3138__delay_3137__delay_3136_reinterpretcast_2560 <= __delay_data_3137__delay_3136_reinterpretcast_2560;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3140__delay_3139_plus_2587 <= __delay_data_3139_plus_2587;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3143__delay_3142__delay_3141__variable_2450 <= __delay_data_3142__delay_3141__variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3156__delay_3155_plus_2592 <= __delay_data_3155_plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3170__delay_3169__delay_3168__variable_2445 <= __delay_data_3169__delay_3168__variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3184__delay_3183__delay_3182_reinterpretcast_2568 <= __delay_data_3183__delay_3182_reinterpretcast_2568;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3186__delay_3185_plus_2613 <= __delay_data_3185_plus_2613;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3189__delay_3188__delay_3187_reinterpretcast_2572 <= __delay_data_3188__delay_3187_reinterpretcast_2572;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3191__delay_3190_plus_2618 <= __delay_data_3190_plus_2618;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3193__delay_3192_plus_2623 <= __delay_data_3192_plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3207__delay_3206__delay_3205_cond_2477 <= __delay_data_3206__delay_3205_cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3227__delay_3226__delay_3225_cond_2489 <= __delay_data_3226__delay_3225_cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3247__delay_3246_plus_2628 <= __delay_data_3246_plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3268__delay_3267_eq_2634 <= __delay_data_3267_eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3300__delay_3299_eq_2637 <= __delay_data_3299_eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3332__delay_3331__delay_3330_cond_2476 <= __delay_data_3331__delay_3330_cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3352__delay_3351__delay_3350_cond_2488 <= __delay_data_3351__delay_3350_cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3372__delay_3371_plus_2597 <= __delay_data_3371_plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3393__delay_3392_eq_2603 <= __delay_data_3392_eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3425__delay_3424_eq_2606 <= __delay_data_3424_eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3144__delay_3143__delay_3142____variable_2450 <= __delay_data_3143__delay_3142__delay_3141__variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3157__delay_3156__delay_3155_plus_2592 <= __delay_data_3156__delay_3155_plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3171__delay_3170__delay_3169____variable_2445 <= __delay_data_3170__delay_3169__delay_3168__variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3194__delay_3193__delay_3192_plus_2623 <= __delay_data_3193__delay_3192_plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3208__delay_3207__delay_3206___cond_2477 <= __delay_data_3207__delay_3206__delay_3205_cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3228__delay_3227__delay_3226___cond_2489 <= __delay_data_3227__delay_3226__delay_3225_cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3248__delay_3247__delay_3246_plus_2628 <= __delay_data_3247__delay_3246_plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3269__delay_3268__delay_3267_eq_2634 <= __delay_data_3268__delay_3267_eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3301__delay_3300__delay_3299_eq_2637 <= __delay_data_3300__delay_3299_eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3333__delay_3332__delay_3331___cond_2476 <= __delay_data_3332__delay_3331__delay_3330_cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3353__delay_3352__delay_3351___cond_2488 <= __delay_data_3352__delay_3351__delay_3350_cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3373__delay_3372__delay_3371_plus_2597 <= __delay_data_3372__delay_3371_plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3394__delay_3393__delay_3392_eq_2603 <= __delay_data_3393__delay_3392_eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3426__delay_3425__delay_3424_eq_2606 <= __delay_data_3425__delay_3424_eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3145__delay_3144__delay_3143____variable_2450 <= __delay_data_3144__delay_3143__delay_3142____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3158__delay_3157__delay_3156___plus_2592 <= __delay_data_3157__delay_3156__delay_3155_plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3172__delay_3171__delay_3170____variable_2445 <= __delay_data_3171__delay_3170__delay_3169____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3195__delay_3194__delay_3193___plus_2623 <= __delay_data_3194__delay_3193__delay_3192_plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3209__delay_3208__delay_3207___cond_2477 <= __delay_data_3208__delay_3207__delay_3206___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3229__delay_3228__delay_3227___cond_2489 <= __delay_data_3228__delay_3227__delay_3226___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3249__delay_3248__delay_3247___plus_2628 <= __delay_data_3248__delay_3247__delay_3246_plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3270__delay_3269__delay_3268__delay_3267_eq_2634 <= __delay_data_3269__delay_3268__delay_3267_eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3302__delay_3301__delay_3300__delay_3299_eq_2637 <= __delay_data_3301__delay_3300__delay_3299_eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3334__delay_3333__delay_3332___cond_2476 <= __delay_data_3333__delay_3332__delay_3331___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3354__delay_3353__delay_3352___cond_2488 <= __delay_data_3353__delay_3352__delay_3351___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3374__delay_3373__delay_3372___plus_2597 <= __delay_data_3373__delay_3372__delay_3371_plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3395__delay_3394__delay_3393__delay_3392_eq_2603 <= __delay_data_3394__delay_3393__delay_3392_eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3427__delay_3426__delay_3425__delay_3424_eq_2606 <= __delay_data_3426__delay_3425__delay_3424_eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3146__delay_3145__delay_3144____variable_2450 <= __delay_data_3145__delay_3144__delay_3143____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3159__delay_3158__delay_3157___plus_2592 <= __delay_data_3158__delay_3157__delay_3156___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3173__delay_3172__delay_3171____variable_2445 <= __delay_data_3172__delay_3171__delay_3170____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3196__delay_3195__delay_3194___plus_2623 <= __delay_data_3195__delay_3194__delay_3193___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3210__delay_3209__delay_3208___cond_2477 <= __delay_data_3209__delay_3208__delay_3207___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3230__delay_3229__delay_3228___cond_2489 <= __delay_data_3229__delay_3228__delay_3227___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3250__delay_3249__delay_3248___plus_2628 <= __delay_data_3249__delay_3248__delay_3247___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3271__delay_3270__delay_3269__delay_3268___eq_2634 <= __delay_data_3270__delay_3269__delay_3268__delay_3267_eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3303__delay_3302__delay_3301__delay_3300___eq_2637 <= __delay_data_3302__delay_3301__delay_3300__delay_3299_eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3335__delay_3334__delay_3333___cond_2476 <= __delay_data_3334__delay_3333__delay_3332___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3355__delay_3354__delay_3353___cond_2488 <= __delay_data_3354__delay_3353__delay_3352___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3375__delay_3374__delay_3373___plus_2597 <= __delay_data_3374__delay_3373__delay_3372___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3396__delay_3395__delay_3394__delay_3393___eq_2603 <= __delay_data_3395__delay_3394__delay_3393__delay_3392_eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3428__delay_3427__delay_3426__delay_3425___eq_2606 <= __delay_data_3427__delay_3426__delay_3425__delay_3424_eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3147__delay_3146__delay_3145____variable_2450 <= __delay_data_3146__delay_3145__delay_3144____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3160__delay_3159__delay_3158___plus_2592 <= __delay_data_3159__delay_3158__delay_3157___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3174__delay_3173__delay_3172____variable_2445 <= __delay_data_3173__delay_3172__delay_3171____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3197__delay_3196__delay_3195___plus_2623 <= __delay_data_3196__delay_3195__delay_3194___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3211__delay_3210__delay_3209___cond_2477 <= __delay_data_3210__delay_3209__delay_3208___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3231__delay_3230__delay_3229___cond_2489 <= __delay_data_3230__delay_3229__delay_3228___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3251__delay_3250__delay_3249___plus_2628 <= __delay_data_3250__delay_3249__delay_3248___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3272__delay_3271__delay_3270__delay_3269___eq_2634 <= __delay_data_3271__delay_3270__delay_3269__delay_3268___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3304__delay_3303__delay_3302__delay_3301___eq_2637 <= __delay_data_3303__delay_3302__delay_3301__delay_3300___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3336__delay_3335__delay_3334___cond_2476 <= __delay_data_3335__delay_3334__delay_3333___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3356__delay_3355__delay_3354___cond_2488 <= __delay_data_3355__delay_3354__delay_3353___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3376__delay_3375__delay_3374___plus_2597 <= __delay_data_3375__delay_3374__delay_3373___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3397__delay_3396__delay_3395__delay_3394___eq_2603 <= __delay_data_3396__delay_3395__delay_3394__delay_3393___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3429__delay_3428__delay_3427__delay_3426___eq_2606 <= __delay_data_3428__delay_3427__delay_3426__delay_3425___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3148__delay_3147__delay_3146____variable_2450 <= __delay_data_3147__delay_3146__delay_3145____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3161__delay_3160__delay_3159___plus_2592 <= __delay_data_3160__delay_3159__delay_3158___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3175__delay_3174__delay_3173____variable_2445 <= __delay_data_3174__delay_3173__delay_3172____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3198__delay_3197__delay_3196___plus_2623 <= __delay_data_3197__delay_3196__delay_3195___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3212__delay_3211__delay_3210___cond_2477 <= __delay_data_3211__delay_3210__delay_3209___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3232__delay_3231__delay_3230___cond_2489 <= __delay_data_3231__delay_3230__delay_3229___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3252__delay_3251__delay_3250___plus_2628 <= __delay_data_3251__delay_3250__delay_3249___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3273__delay_3272__delay_3271__delay_3270___eq_2634 <= __delay_data_3272__delay_3271__delay_3270__delay_3269___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3305__delay_3304__delay_3303__delay_3302___eq_2637 <= __delay_data_3304__delay_3303__delay_3302__delay_3301___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3337__delay_3336__delay_3335___cond_2476 <= __delay_data_3336__delay_3335__delay_3334___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3357__delay_3356__delay_3355___cond_2488 <= __delay_data_3356__delay_3355__delay_3354___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3377__delay_3376__delay_3375___plus_2597 <= __delay_data_3376__delay_3375__delay_3374___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3398__delay_3397__delay_3396__delay_3395___eq_2603 <= __delay_data_3397__delay_3396__delay_3395__delay_3394___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3430__delay_3429__delay_3428__delay_3427___eq_2606 <= __delay_data_3429__delay_3428__delay_3427__delay_3426___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3149__delay_3148__delay_3147____variable_2450 <= __delay_data_3148__delay_3147__delay_3146____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3162__delay_3161__delay_3160___plus_2592 <= __delay_data_3161__delay_3160__delay_3159___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3176__delay_3175__delay_3174____variable_2445 <= __delay_data_3175__delay_3174__delay_3173____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3199__delay_3198__delay_3197___plus_2623 <= __delay_data_3198__delay_3197__delay_3196___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3213__delay_3212__delay_3211___cond_2477 <= __delay_data_3212__delay_3211__delay_3210___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3233__delay_3232__delay_3231___cond_2489 <= __delay_data_3232__delay_3231__delay_3230___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3253__delay_3252__delay_3251___plus_2628 <= __delay_data_3252__delay_3251__delay_3250___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3274__delay_3273__delay_3272__delay_3271___eq_2634 <= __delay_data_3273__delay_3272__delay_3271__delay_3270___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3306__delay_3305__delay_3304__delay_3303___eq_2637 <= __delay_data_3305__delay_3304__delay_3303__delay_3302___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3338__delay_3337__delay_3336___cond_2476 <= __delay_data_3337__delay_3336__delay_3335___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3358__delay_3357__delay_3356___cond_2488 <= __delay_data_3357__delay_3356__delay_3355___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3378__delay_3377__delay_3376___plus_2597 <= __delay_data_3377__delay_3376__delay_3375___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3399__delay_3398__delay_3397__delay_3396___eq_2603 <= __delay_data_3398__delay_3397__delay_3396__delay_3395___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3431__delay_3430__delay_3429__delay_3428___eq_2606 <= __delay_data_3430__delay_3429__delay_3428__delay_3427___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3150__delay_3149__delay_3148____variable_2450 <= __delay_data_3149__delay_3148__delay_3147____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3163__delay_3162__delay_3161___plus_2592 <= __delay_data_3162__delay_3161__delay_3160___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3177__delay_3176__delay_3175____variable_2445 <= __delay_data_3176__delay_3175__delay_3174____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3200__delay_3199__delay_3198___plus_2623 <= __delay_data_3199__delay_3198__delay_3197___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3214__delay_3213__delay_3212___cond_2477 <= __delay_data_3213__delay_3212__delay_3211___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3234__delay_3233__delay_3232___cond_2489 <= __delay_data_3233__delay_3232__delay_3231___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3254__delay_3253__delay_3252___plus_2628 <= __delay_data_3253__delay_3252__delay_3251___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3275__delay_3274__delay_3273__delay_3272___eq_2634 <= __delay_data_3274__delay_3273__delay_3272__delay_3271___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3307__delay_3306__delay_3305__delay_3304___eq_2637 <= __delay_data_3306__delay_3305__delay_3304__delay_3303___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3339__delay_3338__delay_3337___cond_2476 <= __delay_data_3338__delay_3337__delay_3336___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3359__delay_3358__delay_3357___cond_2488 <= __delay_data_3358__delay_3357__delay_3356___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3379__delay_3378__delay_3377___plus_2597 <= __delay_data_3378__delay_3377__delay_3376___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3400__delay_3399__delay_3398__delay_3397___eq_2603 <= __delay_data_3399__delay_3398__delay_3397__delay_3396___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3432__delay_3431__delay_3430__delay_3429___eq_2606 <= __delay_data_3431__delay_3430__delay_3429__delay_3428___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3151__delay_3150__delay_3149____variable_2450 <= __delay_data_3150__delay_3149__delay_3148____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3164__delay_3163__delay_3162___plus_2592 <= __delay_data_3163__delay_3162__delay_3161___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3178__delay_3177__delay_3176____variable_2445 <= __delay_data_3177__delay_3176__delay_3175____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3201__delay_3200__delay_3199___plus_2623 <= __delay_data_3200__delay_3199__delay_3198___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3215__delay_3214__delay_3213___cond_2477 <= __delay_data_3214__delay_3213__delay_3212___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3235__delay_3234__delay_3233___cond_2489 <= __delay_data_3234__delay_3233__delay_3232___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3255__delay_3254__delay_3253___plus_2628 <= __delay_data_3254__delay_3253__delay_3252___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3276__delay_3275__delay_3274__delay_3273___eq_2634 <= __delay_data_3275__delay_3274__delay_3273__delay_3272___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3308__delay_3307__delay_3306__delay_3305___eq_2637 <= __delay_data_3307__delay_3306__delay_3305__delay_3304___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3340__delay_3339__delay_3338___cond_2476 <= __delay_data_3339__delay_3338__delay_3337___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3360__delay_3359__delay_3358___cond_2488 <= __delay_data_3359__delay_3358__delay_3357___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3380__delay_3379__delay_3378___plus_2597 <= __delay_data_3379__delay_3378__delay_3377___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3401__delay_3400__delay_3399__delay_3398___eq_2603 <= __delay_data_3400__delay_3399__delay_3398__delay_3397___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3433__delay_3432__delay_3431__delay_3430___eq_2606 <= __delay_data_3432__delay_3431__delay_3430__delay_3429___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3152__delay_3151__delay_3150____variable_2450 <= __delay_data_3151__delay_3150__delay_3149____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3165__delay_3164__delay_3163___plus_2592 <= __delay_data_3164__delay_3163__delay_3162___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3179__delay_3178__delay_3177____variable_2445 <= __delay_data_3178__delay_3177__delay_3176____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3202__delay_3201__delay_3200___plus_2623 <= __delay_data_3201__delay_3200__delay_3199___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3216__delay_3215__delay_3214___cond_2477 <= __delay_data_3215__delay_3214__delay_3213___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3236__delay_3235__delay_3234___cond_2489 <= __delay_data_3235__delay_3234__delay_3233___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3256__delay_3255__delay_3254___plus_2628 <= __delay_data_3255__delay_3254__delay_3253___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3277__delay_3276__delay_3275__delay_3274___eq_2634 <= __delay_data_3276__delay_3275__delay_3274__delay_3273___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3309__delay_3308__delay_3307__delay_3306___eq_2637 <= __delay_data_3308__delay_3307__delay_3306__delay_3305___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3341__delay_3340__delay_3339___cond_2476 <= __delay_data_3340__delay_3339__delay_3338___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3361__delay_3360__delay_3359___cond_2488 <= __delay_data_3360__delay_3359__delay_3358___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3381__delay_3380__delay_3379___plus_2597 <= __delay_data_3380__delay_3379__delay_3378___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3402__delay_3401__delay_3400__delay_3399___eq_2603 <= __delay_data_3401__delay_3400__delay_3399__delay_3398___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3434__delay_3433__delay_3432__delay_3431___eq_2606 <= __delay_data_3433__delay_3432__delay_3431__delay_3430___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3153__delay_3152__delay_3151____variable_2450 <= __delay_data_3152__delay_3151__delay_3150____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3166__delay_3165__delay_3164___plus_2592 <= __delay_data_3165__delay_3164__delay_3163___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3180__delay_3179__delay_3178____variable_2445 <= __delay_data_3179__delay_3178__delay_3177____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3203__delay_3202__delay_3201___plus_2623 <= __delay_data_3202__delay_3201__delay_3200___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3217__delay_3216__delay_3215___cond_2477 <= __delay_data_3216__delay_3215__delay_3214___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3237__delay_3236__delay_3235___cond_2489 <= __delay_data_3236__delay_3235__delay_3234___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3257__delay_3256__delay_3255___plus_2628 <= __delay_data_3256__delay_3255__delay_3254___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3278__delay_3277__delay_3276__delay_3275___eq_2634 <= __delay_data_3277__delay_3276__delay_3275__delay_3274___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3310__delay_3309__delay_3308__delay_3307___eq_2637 <= __delay_data_3309__delay_3308__delay_3307__delay_3306___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3342__delay_3341__delay_3340___cond_2476 <= __delay_data_3341__delay_3340__delay_3339___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3362__delay_3361__delay_3360___cond_2488 <= __delay_data_3361__delay_3360__delay_3359___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3382__delay_3381__delay_3380___plus_2597 <= __delay_data_3381__delay_3380__delay_3379___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3403__delay_3402__delay_3401__delay_3400___eq_2603 <= __delay_data_3402__delay_3401__delay_3400__delay_3399___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3435__delay_3434__delay_3433__delay_3432___eq_2606 <= __delay_data_3434__delay_3433__delay_3432__delay_3431___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3154__delay_3153__delay_3152____variable_2450 <= __delay_data_3153__delay_3152__delay_3151____variable_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3167__delay_3166__delay_3165___plus_2592 <= __delay_data_3166__delay_3165__delay_3164___plus_2592;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3181__delay_3180__delay_3179____variable_2445 <= __delay_data_3180__delay_3179__delay_3178____variable_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3204__delay_3203__delay_3202___plus_2623 <= __delay_data_3203__delay_3202__delay_3201___plus_2623;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3218__delay_3217__delay_3216___cond_2477 <= __delay_data_3217__delay_3216__delay_3215___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3238__delay_3237__delay_3236___cond_2489 <= __delay_data_3237__delay_3236__delay_3235___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3258__delay_3257__delay_3256___plus_2628 <= __delay_data_3257__delay_3256__delay_3255___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3279__delay_3278__delay_3277__delay_3276___eq_2634 <= __delay_data_3278__delay_3277__delay_3276__delay_3275___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3311__delay_3310__delay_3309__delay_3308___eq_2637 <= __delay_data_3310__delay_3309__delay_3308__delay_3307___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3343__delay_3342__delay_3341___cond_2476 <= __delay_data_3342__delay_3341__delay_3340___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3363__delay_3362__delay_3361___cond_2488 <= __delay_data_3362__delay_3361__delay_3360___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3383__delay_3382__delay_3381___plus_2597 <= __delay_data_3382__delay_3381__delay_3380___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3404__delay_3403__delay_3402__delay_3401___eq_2603 <= __delay_data_3403__delay_3402__delay_3401__delay_3400___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3436__delay_3435__delay_3434__delay_3433___eq_2606 <= __delay_data_3435__delay_3434__delay_3433__delay_3432___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3219__delay_3218__delay_3217___cond_2477 <= __delay_data_3218__delay_3217__delay_3216___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3239__delay_3238__delay_3237___cond_2489 <= __delay_data_3238__delay_3237__delay_3236___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3259__delay_3258__delay_3257___plus_2628 <= __delay_data_3258__delay_3257__delay_3256___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3280__delay_3279__delay_3278__delay_3277___eq_2634 <= __delay_data_3279__delay_3278__delay_3277__delay_3276___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3312__delay_3311__delay_3310__delay_3309___eq_2637 <= __delay_data_3311__delay_3310__delay_3309__delay_3308___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3344__delay_3343__delay_3342___cond_2476 <= __delay_data_3343__delay_3342__delay_3341___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3364__delay_3363__delay_3362___cond_2488 <= __delay_data_3363__delay_3362__delay_3361___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3384__delay_3383__delay_3382___plus_2597 <= __delay_data_3383__delay_3382__delay_3381___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3405__delay_3404__delay_3403__delay_3402___eq_2603 <= __delay_data_3404__delay_3403__delay_3402__delay_3401___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3437__delay_3436__delay_3435__delay_3434___eq_2606 <= __delay_data_3436__delay_3435__delay_3434__delay_3433___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3220__delay_3219__delay_3218___cond_2477 <= __delay_data_3219__delay_3218__delay_3217___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3240__delay_3239__delay_3238___cond_2489 <= __delay_data_3239__delay_3238__delay_3237___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3260__delay_3259__delay_3258___plus_2628 <= __delay_data_3259__delay_3258__delay_3257___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3281__delay_3280__delay_3279__delay_3278___eq_2634 <= __delay_data_3280__delay_3279__delay_3278__delay_3277___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3313__delay_3312__delay_3311__delay_3310___eq_2637 <= __delay_data_3312__delay_3311__delay_3310__delay_3309___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3345__delay_3344__delay_3343___cond_2476 <= __delay_data_3344__delay_3343__delay_3342___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3365__delay_3364__delay_3363___cond_2488 <= __delay_data_3364__delay_3363__delay_3362___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3385__delay_3384__delay_3383___plus_2597 <= __delay_data_3384__delay_3383__delay_3382___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3406__delay_3405__delay_3404__delay_3403___eq_2603 <= __delay_data_3405__delay_3404__delay_3403__delay_3402___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3438__delay_3437__delay_3436__delay_3435___eq_2606 <= __delay_data_3437__delay_3436__delay_3435__delay_3434___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3221__delay_3220__delay_3219___cond_2477 <= __delay_data_3220__delay_3219__delay_3218___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3241__delay_3240__delay_3239___cond_2489 <= __delay_data_3240__delay_3239__delay_3238___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3261__delay_3260__delay_3259___plus_2628 <= __delay_data_3260__delay_3259__delay_3258___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3282__delay_3281__delay_3280__delay_3279___eq_2634 <= __delay_data_3281__delay_3280__delay_3279__delay_3278___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3314__delay_3313__delay_3312__delay_3311___eq_2637 <= __delay_data_3313__delay_3312__delay_3311__delay_3310___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3346__delay_3345__delay_3344___cond_2476 <= __delay_data_3345__delay_3344__delay_3343___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3366__delay_3365__delay_3364___cond_2488 <= __delay_data_3365__delay_3364__delay_3363___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3386__delay_3385__delay_3384___plus_2597 <= __delay_data_3385__delay_3384__delay_3383___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3407__delay_3406__delay_3405__delay_3404___eq_2603 <= __delay_data_3406__delay_3405__delay_3404__delay_3403___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3439__delay_3438__delay_3437__delay_3436___eq_2606 <= __delay_data_3438__delay_3437__delay_3436__delay_3435___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3222__delay_3221__delay_3220___cond_2477 <= __delay_data_3221__delay_3220__delay_3219___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3242__delay_3241__delay_3240___cond_2489 <= __delay_data_3241__delay_3240__delay_3239___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3262__delay_3261__delay_3260___plus_2628 <= __delay_data_3261__delay_3260__delay_3259___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3283__delay_3282__delay_3281__delay_3280___eq_2634 <= __delay_data_3282__delay_3281__delay_3280__delay_3279___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3315__delay_3314__delay_3313__delay_3312___eq_2637 <= __delay_data_3314__delay_3313__delay_3312__delay_3311___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3347__delay_3346__delay_3345___cond_2476 <= __delay_data_3346__delay_3345__delay_3344___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3367__delay_3366__delay_3365___cond_2488 <= __delay_data_3366__delay_3365__delay_3364___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3387__delay_3386__delay_3385___plus_2597 <= __delay_data_3386__delay_3385__delay_3384___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3408__delay_3407__delay_3406__delay_3405___eq_2603 <= __delay_data_3407__delay_3406__delay_3405__delay_3404___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3440__delay_3439__delay_3438__delay_3437___eq_2606 <= __delay_data_3439__delay_3438__delay_3437__delay_3436___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3223__delay_3222__delay_3221___cond_2477 <= __delay_data_3222__delay_3221__delay_3220___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3243__delay_3242__delay_3241___cond_2489 <= __delay_data_3242__delay_3241__delay_3240___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3263__delay_3262__delay_3261___plus_2628 <= __delay_data_3262__delay_3261__delay_3260___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3284__delay_3283__delay_3282__delay_3281___eq_2634 <= __delay_data_3283__delay_3282__delay_3281__delay_3280___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3316__delay_3315__delay_3314__delay_3313___eq_2637 <= __delay_data_3315__delay_3314__delay_3313__delay_3312___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3348__delay_3347__delay_3346___cond_2476 <= __delay_data_3347__delay_3346__delay_3345___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3368__delay_3367__delay_3366___cond_2488 <= __delay_data_3367__delay_3366__delay_3365___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3388__delay_3387__delay_3386___plus_2597 <= __delay_data_3387__delay_3386__delay_3385___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3409__delay_3408__delay_3407__delay_3406___eq_2603 <= __delay_data_3408__delay_3407__delay_3406__delay_3405___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3441__delay_3440__delay_3439__delay_3438___eq_2606 <= __delay_data_3440__delay_3439__delay_3438__delay_3437___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3224__delay_3223__delay_3222___cond_2477 <= __delay_data_3223__delay_3222__delay_3221___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3244__delay_3243__delay_3242___cond_2489 <= __delay_data_3243__delay_3242__delay_3241___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3264__delay_3263__delay_3262___plus_2628 <= __delay_data_3263__delay_3262__delay_3261___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3285__delay_3284__delay_3283__delay_3282___eq_2634 <= __delay_data_3284__delay_3283__delay_3282__delay_3281___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3317__delay_3316__delay_3315__delay_3314___eq_2637 <= __delay_data_3316__delay_3315__delay_3314__delay_3313___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3349__delay_3348__delay_3347___cond_2476 <= __delay_data_3348__delay_3347__delay_3346___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3369__delay_3368__delay_3367___cond_2488 <= __delay_data_3368__delay_3367__delay_3366___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3389__delay_3388__delay_3387___plus_2597 <= __delay_data_3388__delay_3387__delay_3386___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3410__delay_3409__delay_3408__delay_3407___eq_2603 <= __delay_data_3409__delay_3408__delay_3407__delay_3406___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3442__delay_3441__delay_3440__delay_3439___eq_2606 <= __delay_data_3441__delay_3440__delay_3439__delay_3438___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2595 <= __substreamoutput_data_2593 + __delay_data_3349__delay_3348__delay_3347___cond_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _plus_data_2626 <= __substreamoutput_data_2624 + __delay_data_3224__delay_3223__delay_3222___cond_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3245__delay_3244__delay_3243___cond_2489 <= __delay_data_3244__delay_3243__delay_3242___cond_2489;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3265__delay_3264__delay_3263___plus_2628 <= __delay_data_3264__delay_3263__delay_3262___plus_2628;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3286__delay_3285__delay_3284__delay_3283___eq_2634 <= __delay_data_3285__delay_3284__delay_3283__delay_3282___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3318__delay_3317__delay_3316__delay_3315___eq_2637 <= __delay_data_3317__delay_3316__delay_3315__delay_3314___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3370__delay_3369__delay_3368___cond_2488 <= __delay_data_3369__delay_3368__delay_3367___cond_2488;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3390__delay_3389__delay_3388___plus_2597 <= __delay_data_3389__delay_3388__delay_3387___plus_2597;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3411__delay_3410__delay_3409__delay_3408___eq_2603 <= __delay_data_3410__delay_3409__delay_3408__delay_3407___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3443__delay_3442__delay_3441__delay_3440___eq_2606 <= __delay_data_3442__delay_3441__delay_3440__delay_3439___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3455__substreamoutput_2594 <= __substreamoutput_data_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3287__delay_3286__delay_3285__delay_3284___eq_2634 <= __delay_data_3286__delay_3285__delay_3284__delay_3283___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3319__delay_3318__delay_3317__delay_3316___eq_2637 <= __delay_data_3318__delay_3317__delay_3316__delay_3315___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3412__delay_3411__delay_3410__delay_3409___eq_2603 <= __delay_data_3411__delay_3410__delay_3409__delay_3408___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3444__delay_3443__delay_3442__delay_3441___eq_2606 <= __delay_data_3443__delay_3442__delay_3441__delay_3440___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3456__delay_3455__substreamoutput_2594 <= __delay_data_3455__substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3288__delay_3287__delay_3286__delay_3285___eq_2634 <= __delay_data_3287__delay_3286__delay_3285__delay_3284___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3320__delay_3319__delay_3318__delay_3317___eq_2637 <= __delay_data_3319__delay_3318__delay_3317__delay_3316___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3413__delay_3412__delay_3411__delay_3410___eq_2603 <= __delay_data_3412__delay_3411__delay_3410__delay_3409___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3445__delay_3444__delay_3443__delay_3442___eq_2606 <= __delay_data_3444__delay_3443__delay_3442__delay_3441___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3457__delay_3456____substreamoutput_2594 <= __delay_data_3456__delay_3455__substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3289__delay_3288__delay_3287__delay_3286___eq_2634 <= __delay_data_3288__delay_3287__delay_3286__delay_3285___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3321__delay_3320__delay_3319__delay_3318___eq_2637 <= __delay_data_3320__delay_3319__delay_3318__delay_3317___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3414__delay_3413__delay_3412__delay_3411___eq_2603 <= __delay_data_3413__delay_3412__delay_3411__delay_3410___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3446__delay_3445__delay_3444__delay_3443___eq_2606 <= __delay_data_3445__delay_3444__delay_3443__delay_3442___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3458__delay_3457____substreamoutput_2594 <= __delay_data_3457__delay_3456____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3290__delay_3289__delay_3288__delay_3287___eq_2634 <= __delay_data_3289__delay_3288__delay_3287__delay_3286___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3322__delay_3321__delay_3320__delay_3319___eq_2637 <= __delay_data_3321__delay_3320__delay_3319__delay_3318___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3415__delay_3414__delay_3413__delay_3412___eq_2603 <= __delay_data_3414__delay_3413__delay_3412__delay_3411___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3447__delay_3446__delay_3445__delay_3444___eq_2606 <= __delay_data_3446__delay_3445__delay_3444__delay_3443___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3459__delay_3458____substreamoutput_2594 <= __delay_data_3458__delay_3457____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3291__delay_3290__delay_3289__delay_3288___eq_2634 <= __delay_data_3290__delay_3289__delay_3288__delay_3287___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3323__delay_3322__delay_3321__delay_3320___eq_2637 <= __delay_data_3322__delay_3321__delay_3320__delay_3319___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3416__delay_3415__delay_3414__delay_3413___eq_2603 <= __delay_data_3415__delay_3414__delay_3413__delay_3412___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3448__delay_3447__delay_3446__delay_3445___eq_2606 <= __delay_data_3447__delay_3446__delay_3445__delay_3444___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3460__delay_3459____substreamoutput_2594 <= __delay_data_3459__delay_3458____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3292__delay_3291__delay_3290__delay_3289___eq_2634 <= __delay_data_3291__delay_3290__delay_3289__delay_3288___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3324__delay_3323__delay_3322__delay_3321___eq_2637 <= __delay_data_3323__delay_3322__delay_3321__delay_3320___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3417__delay_3416__delay_3415__delay_3414___eq_2603 <= __delay_data_3416__delay_3415__delay_3414__delay_3413___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3449__delay_3448__delay_3447__delay_3446___eq_2606 <= __delay_data_3448__delay_3447__delay_3446__delay_3445___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3461__delay_3460____substreamoutput_2594 <= __delay_data_3460__delay_3459____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3293__delay_3292__delay_3291__delay_3290___eq_2634 <= __delay_data_3292__delay_3291__delay_3290__delay_3289___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3325__delay_3324__delay_3323__delay_3322___eq_2637 <= __delay_data_3324__delay_3323__delay_3322__delay_3321___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3418__delay_3417__delay_3416__delay_3415___eq_2603 <= __delay_data_3417__delay_3416__delay_3415__delay_3414___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3450__delay_3449__delay_3448__delay_3447___eq_2606 <= __delay_data_3449__delay_3448__delay_3447__delay_3446___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3462__delay_3461____substreamoutput_2594 <= __delay_data_3461__delay_3460____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3294__delay_3293__delay_3292__delay_3291___eq_2634 <= __delay_data_3293__delay_3292__delay_3291__delay_3290___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3326__delay_3325__delay_3324__delay_3323___eq_2637 <= __delay_data_3325__delay_3324__delay_3323__delay_3322___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3419__delay_3418__delay_3417__delay_3416___eq_2603 <= __delay_data_3418__delay_3417__delay_3416__delay_3415___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3451__delay_3450__delay_3449__delay_3448___eq_2606 <= __delay_data_3450__delay_3449__delay_3448__delay_3447___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3463__delay_3462____substreamoutput_2594 <= __delay_data_3462__delay_3461____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3295__delay_3294__delay_3293__delay_3292___eq_2634 <= __delay_data_3294__delay_3293__delay_3292__delay_3291___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3327__delay_3326__delay_3325__delay_3324___eq_2637 <= __delay_data_3326__delay_3325__delay_3324__delay_3323___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3420__delay_3419__delay_3418__delay_3417___eq_2603 <= __delay_data_3419__delay_3418__delay_3417__delay_3416___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3452__delay_3451__delay_3450__delay_3449___eq_2606 <= __delay_data_3451__delay_3450__delay_3449__delay_3448___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3464__delay_3463____substreamoutput_2594 <= __delay_data_3463__delay_3462____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _greaterthan_data_2600 <= __substreamoutput_data_2598 > 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _greaterthan_data_2631 <= __substreamoutput_data_2629 > 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3266__substreamoutput_2629 <= __substreamoutput_data_2629;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3296__delay_3295__delay_3294__delay_3293___eq_2634 <= __delay_data_3295__delay_3294__delay_3293__delay_3292___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3328__delay_3327__delay_3326__delay_3325___eq_2637 <= __delay_data_3327__delay_3326__delay_3325__delay_3324___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3391__substreamoutput_2598 <= __substreamoutput_data_2598;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3421__delay_3420__delay_3419__delay_3418___eq_2603 <= __delay_data_3420__delay_3419__delay_3418__delay_3417___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3453__delay_3452__delay_3451__delay_3450___eq_2606 <= __delay_data_3452__delay_3451__delay_3450__delay_3449___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3465__delay_3464____substreamoutput_2594 <= __delay_data_3464__delay_3463____substreamoutput_2594;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _cond_data_2602 <= (_greaterthan_data_2600)? __delay_data_3391__substreamoutput_2598 : 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _cond_data_2633 <= (_greaterthan_data_2631)? __delay_data_3266__substreamoutput_2629 : 1'sd0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3297__delay_3296__delay_3295__delay_3294___eq_2634 <= __delay_data_3296__delay_3295__delay_3294__delay_3293___eq_2634;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3298__delay_3266__substreamoutput_2629 <= __delay_data_3266__substreamoutput_2629;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3329__delay_3328__delay_3327__delay_3326___eq_2637 <= __delay_data_3328__delay_3327__delay_3326__delay_3325___eq_2637;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3422__delay_3421__delay_3420__delay_3419___eq_2603 <= __delay_data_3421__delay_3420__delay_3419__delay_3418___eq_2603;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3423__delay_3391__substreamoutput_2598 <= __delay_data_3391__substreamoutput_2598;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3454__delay_3453__delay_3452__delay_3451___eq_2606 <= __delay_data_3453__delay_3452__delay_3451__delay_3450___eq_2606;
      end 
      if(_stream_matmul_16_stream_oready) begin
        __delay_data_3466__delay_3465____substreamoutput_2594 <= __delay_data_3465__delay_3464____substreamoutput_2594;
      end 
      if(_set_flag_2207) begin
        _stream_matmul_16_parameter_0_next_parameter_data <= cparam_matmul_16_stream_reduce_size;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2445 <= _stream_matmul_16_parameter_0_next_parameter_data;
      end 
      if(_set_flag_2208) begin
        _stream_matmul_16_parameter_1_next_parameter_data <= matmul_16_col_select;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2446 <= _stream_matmul_16_parameter_1_next_parameter_data;
      end 
      if(_set_flag_2209) begin
        _stream_matmul_16_parameter_2_next_parameter_data <= matmul_16_row_select_buf;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2447 <= _stream_matmul_16_parameter_2_next_parameter_data;
      end 
      if(_set_flag_2210) begin
        _stream_matmul_16_parameter_3_next_parameter_data <= matmul_16_stream_pad_masks;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2448 <= _stream_matmul_16_parameter_3_next_parameter_data;
      end 
      if(_set_flag_2211) begin
        _stream_matmul_16_parameter_4_next_parameter_data <= cparam_matmul_16_stream_omit_mask;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2449 <= _stream_matmul_16_parameter_4_next_parameter_data;
      end 
      if(_set_flag_2212) begin
        _stream_matmul_16_parameter_6_next_parameter_data <= cparam_matmul_16_bias_scala;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2466 <= _stream_matmul_16_parameter_6_next_parameter_data;
      end 
      if(_set_flag_2213) begin
        _stream_matmul_16_source_7_source_mode <= 5'b10;
        _stream_matmul_16_source_7_source_offset <= (cparam_matmul_16_bias_num == 1)? 0 : matmul_16_och_count_buf;
      end 
      if(_set_flag_2213) begin
        _source_stream_matmul_16_source_7_pat_size_0 <= cparam_matmul_16_stream_reduce_size;
        _source_stream_matmul_16_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_2213) begin
        _source_stream_matmul_16_source_7_pat_size_1 <= matmul_16_next_stream_num_ops;
        _source_stream_matmul_16_source_7_pat_stride_1 <= (cparam_matmul_16_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_2213) begin
        _source_stream_matmul_16_source_7_pat_size_2 <= 1;
        _source_stream_matmul_16_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_2213) begin
        _source_stream_matmul_16_source_7_pat_size_3 <= 1;
        _source_stream_matmul_16_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_2213) begin
        _stream_matmul_16_source_7_source_sel <= 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_7_source_offset_buf <= _stream_matmul_16_source_7_source_offset;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_count_0 <= _source_stream_matmul_16_source_7_pat_size_0 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_count_1 <= _source_stream_matmul_16_source_7_pat_size_1 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_count_2 <= _source_stream_matmul_16_source_7_pat_size_2 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_count_3 <= _source_stream_matmul_16_source_7_pat_size_3 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_size_buf_0 <= _source_stream_matmul_16_source_7_pat_size_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_size_buf_1 <= _source_stream_matmul_16_source_7_pat_size_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_size_buf_2 <= _source_stream_matmul_16_source_7_pat_size_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_size_buf_3 <= _source_stream_matmul_16_source_7_pat_size_3;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_stride_buf_0 <= _source_stream_matmul_16_source_7_pat_stride_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_stride_buf_1 <= _source_stream_matmul_16_source_7_pat_stride_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_stride_buf_2 <= _source_stream_matmul_16_source_7_pat_stride_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_stride_buf_3 <= _source_stream_matmul_16_source_7_pat_stride_3;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_source_busy && _stream_matmul_16_is_root) begin
        __variable_wdata_2467 <= _stream_matmul_16_source_7_source_ram_rdata;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_7_idle <= 0;
        _stream_matmul_16_source_7_source_ram_raddr <= _stream_matmul_16_source_7_source_pat_all_offset;
        _stream_matmul_16_source_7_source_ram_renable <= 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_0 <= _source_stream_matmul_16_source_7_pat_cur_offset_0 + _source_stream_matmul_16_source_7_pat_stride_buf_0;
        _source_stream_matmul_16_source_7_pat_count_0 <= _source_stream_matmul_16_source_7_pat_count_0 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_16_source_7_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_0 <= 0;
        _source_stream_matmul_16_source_7_pat_count_0 <= _source_stream_matmul_16_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_16_source_7_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_1 <= _source_stream_matmul_16_source_7_pat_cur_offset_1 + _source_stream_matmul_16_source_7_pat_stride_buf_1;
        _source_stream_matmul_16_source_7_pat_count_1 <= _source_stream_matmul_16_source_7_pat_count_1 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_16_source_7_pat_count_0 == 0) && (_source_stream_matmul_16_source_7_pat_count_1 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_1 <= 0;
        _source_stream_matmul_16_source_7_pat_count_1 <= _source_stream_matmul_16_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_16_source_7_pat_count_0 == 0) && (_source_stream_matmul_16_source_7_pat_count_1 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_2 <= _source_stream_matmul_16_source_7_pat_cur_offset_2 + _source_stream_matmul_16_source_7_pat_stride_buf_2;
        _source_stream_matmul_16_source_7_pat_count_2 <= _source_stream_matmul_16_source_7_pat_count_2 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_16_source_7_pat_count_0 == 0) && (_source_stream_matmul_16_source_7_pat_count_1 == 0)) && (_source_stream_matmul_16_source_7_pat_count_2 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_2 <= 0;
        _source_stream_matmul_16_source_7_pat_count_2 <= _source_stream_matmul_16_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_16_source_7_pat_count_0 == 0) && (_source_stream_matmul_16_source_7_pat_count_1 == 0) && (_source_stream_matmul_16_source_7_pat_count_2 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_3 <= _source_stream_matmul_16_source_7_pat_cur_offset_3 + _source_stream_matmul_16_source_7_pat_stride_buf_3;
        _source_stream_matmul_16_source_7_pat_count_3 <= _source_stream_matmul_16_source_7_pat_count_3 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_16_source_7_pat_count_0 == 0) && (_source_stream_matmul_16_source_7_pat_count_1 == 0) && (_source_stream_matmul_16_source_7_pat_count_2 == 0)) && (_source_stream_matmul_16_source_7_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_7_pat_cur_offset_3 <= 0;
        _source_stream_matmul_16_source_7_pat_count_3 <= _source_stream_matmul_16_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 1) && _stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_7_source_ram_renable <= 0;
        _stream_matmul_16_source_7_idle <= 1;
      end 
      if((_stream_matmul_16_source_7_source_pat_fsm_0 == 2) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_7_source_ram_renable <= 0;
        _stream_matmul_16_source_7_idle <= 1;
      end 
      if(_set_flag_2216) begin
        _stream_matmul_16_parameter_8_next_parameter_data <= cparam_matmul_16_scale_scala;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2478 <= _stream_matmul_16_parameter_8_next_parameter_data;
      end 
      if(_set_flag_2217) begin
        _stream_matmul_16_source_9_source_mode <= 5'b10;
        _stream_matmul_16_source_9_source_offset <= (cparam_matmul_16_scale_num == 1)? 0 : matmul_16_och_count_buf;
      end 
      if(_set_flag_2217) begin
        _source_stream_matmul_16_source_9_pat_size_0 <= cparam_matmul_16_stream_reduce_size;
        _source_stream_matmul_16_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_2217) begin
        _source_stream_matmul_16_source_9_pat_size_1 <= matmul_16_next_stream_num_ops;
        _source_stream_matmul_16_source_9_pat_stride_1 <= (cparam_matmul_16_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_2217) begin
        _source_stream_matmul_16_source_9_pat_size_2 <= 1;
        _source_stream_matmul_16_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_2217) begin
        _source_stream_matmul_16_source_9_pat_size_3 <= 1;
        _source_stream_matmul_16_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_2217) begin
        _stream_matmul_16_source_9_source_sel <= 2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_9_source_offset_buf <= _stream_matmul_16_source_9_source_offset;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_count_0 <= _source_stream_matmul_16_source_9_pat_size_0 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_count_1 <= _source_stream_matmul_16_source_9_pat_size_1 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_count_2 <= _source_stream_matmul_16_source_9_pat_size_2 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_count_3 <= _source_stream_matmul_16_source_9_pat_size_3 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_size_buf_0 <= _source_stream_matmul_16_source_9_pat_size_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_size_buf_1 <= _source_stream_matmul_16_source_9_pat_size_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_size_buf_2 <= _source_stream_matmul_16_source_9_pat_size_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_size_buf_3 <= _source_stream_matmul_16_source_9_pat_size_3;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_stride_buf_0 <= _source_stream_matmul_16_source_9_pat_stride_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_stride_buf_1 <= _source_stream_matmul_16_source_9_pat_stride_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_stride_buf_2 <= _source_stream_matmul_16_source_9_pat_stride_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_stride_buf_3 <= _source_stream_matmul_16_source_9_pat_stride_3;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_source_busy && _stream_matmul_16_is_root) begin
        __variable_wdata_2479 <= _stream_matmul_16_source_9_source_ram_rdata;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_9_idle <= 0;
        _stream_matmul_16_source_9_source_ram_raddr <= _stream_matmul_16_source_9_source_pat_all_offset;
        _stream_matmul_16_source_9_source_ram_renable <= 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_0 <= _source_stream_matmul_16_source_9_pat_cur_offset_0 + _source_stream_matmul_16_source_9_pat_stride_buf_0;
        _source_stream_matmul_16_source_9_pat_count_0 <= _source_stream_matmul_16_source_9_pat_count_0 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_16_source_9_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_0 <= 0;
        _source_stream_matmul_16_source_9_pat_count_0 <= _source_stream_matmul_16_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_16_source_9_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_1 <= _source_stream_matmul_16_source_9_pat_cur_offset_1 + _source_stream_matmul_16_source_9_pat_stride_buf_1;
        _source_stream_matmul_16_source_9_pat_count_1 <= _source_stream_matmul_16_source_9_pat_count_1 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_16_source_9_pat_count_0 == 0) && (_source_stream_matmul_16_source_9_pat_count_1 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_1 <= 0;
        _source_stream_matmul_16_source_9_pat_count_1 <= _source_stream_matmul_16_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_16_source_9_pat_count_0 == 0) && (_source_stream_matmul_16_source_9_pat_count_1 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_2 <= _source_stream_matmul_16_source_9_pat_cur_offset_2 + _source_stream_matmul_16_source_9_pat_stride_buf_2;
        _source_stream_matmul_16_source_9_pat_count_2 <= _source_stream_matmul_16_source_9_pat_count_2 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_16_source_9_pat_count_0 == 0) && (_source_stream_matmul_16_source_9_pat_count_1 == 0)) && (_source_stream_matmul_16_source_9_pat_count_2 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_2 <= 0;
        _source_stream_matmul_16_source_9_pat_count_2 <= _source_stream_matmul_16_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_16_source_9_pat_count_0 == 0) && (_source_stream_matmul_16_source_9_pat_count_1 == 0) && (_source_stream_matmul_16_source_9_pat_count_2 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_3 <= _source_stream_matmul_16_source_9_pat_cur_offset_3 + _source_stream_matmul_16_source_9_pat_stride_buf_3;
        _source_stream_matmul_16_source_9_pat_count_3 <= _source_stream_matmul_16_source_9_pat_count_3 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_16_source_9_pat_count_0 == 0) && (_source_stream_matmul_16_source_9_pat_count_1 == 0) && (_source_stream_matmul_16_source_9_pat_count_2 == 0)) && (_source_stream_matmul_16_source_9_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_9_pat_cur_offset_3 <= 0;
        _source_stream_matmul_16_source_9_pat_count_3 <= _source_stream_matmul_16_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 1) && _stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_9_source_ram_renable <= 0;
        _stream_matmul_16_source_9_idle <= 1;
      end 
      if((_stream_matmul_16_source_9_source_pat_fsm_1 == 2) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_9_source_ram_renable <= 0;
        _stream_matmul_16_source_9_idle <= 1;
      end 
      if(_set_flag_2220) begin
        _stream_matmul_16_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2490 <= _stream_matmul_16_parameter_10_next_parameter_data;
      end 
      if(_set_flag_2221) begin
        _stream_matmul_16_source_11_source_mode <= 5'b0;
        _stream_matmul_16_source_11_source_empty_data <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready && !(|(_stream_matmul_16_source_11_source_mode & 5'b0))) begin
        _stream_matmul_16_source_11_idle <= 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready && !(|(_stream_matmul_16_source_11_source_mode & 5'b0)) && _stream_matmul_16_is_root) begin
        __variable_wdata_2491 <= _stream_matmul_16_source_11_source_empty_data;
      end 
      if(_set_flag_2222) begin
        _stream_matmul_16_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2502 <= _stream_matmul_16_parameter_12_next_parameter_data;
      end 
      if(_set_flag_2223) begin
        _stream_matmul_16_source_13_source_mode <= 5'b0;
        _stream_matmul_16_source_13_source_empty_data <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready && !(|(_stream_matmul_16_source_13_source_mode & 5'b0))) begin
        _stream_matmul_16_source_13_idle <= 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready && !(|(_stream_matmul_16_source_13_source_mode & 5'b0)) && _stream_matmul_16_is_root) begin
        __variable_wdata_2503 <= _stream_matmul_16_source_13_source_empty_data;
      end 
      if(_set_flag_2224) begin
        _stream_matmul_16_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2514 <= _stream_matmul_16_parameter_14_next_parameter_data;
      end 
      if(_set_flag_2225) begin
        _stream_matmul_16_source_15_source_mode <= 5'b0;
        _stream_matmul_16_source_15_source_empty_data <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready && !(|(_stream_matmul_16_source_15_source_mode & 5'b0))) begin
        _stream_matmul_16_source_15_idle <= 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready && !(|(_stream_matmul_16_source_15_source_mode & 5'b0)) && _stream_matmul_16_is_root) begin
        __variable_wdata_2515 <= _stream_matmul_16_source_15_source_empty_data;
      end 
      if(_set_flag_2226) begin
        _stream_matmul_16_parameter_16_next_parameter_data <= cparam_matmul_16_cshamt_mul_value;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2526 <= _stream_matmul_16_parameter_16_next_parameter_data;
      end 
      if(_set_flag_2227) begin
        _stream_matmul_16_parameter_17_next_parameter_data <= cparam_matmul_16_cshamt_sum_value;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2527 <= _stream_matmul_16_parameter_17_next_parameter_data;
      end 
      if(_set_flag_2228) begin
        _stream_matmul_16_parameter_18_next_parameter_data <= cparam_matmul_16_cshamt_out_value;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2528 <= _stream_matmul_16_parameter_18_next_parameter_data;
      end 
      if(_set_flag_2229) begin
        _stream_matmul_16_parameter_19_next_parameter_data <= cparam_matmul_16_act_func_index;
      end 
      if(_stream_matmul_16_source_start) begin
        __variable_wdata_2529 <= _stream_matmul_16_parameter_19_next_parameter_data;
      end 
      if(_set_flag_2230) begin
        _stream_matmul_16_source_20_source_mode <= 5'b10;
        _stream_matmul_16_source_20_source_offset <= matmul_16_stream_act_local_0 + matmul_16_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_2230) begin
        _source_stream_matmul_16_source_20_pat_size_0 <= cparam_matmul_16_stream_reduce_size;
        _source_stream_matmul_16_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_2230) begin
        _source_stream_matmul_16_source_20_pat_size_1 <= matmul_16_next_stream_num_ops;
        _source_stream_matmul_16_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_2230) begin
        _source_stream_matmul_16_source_20_pat_size_2 <= 1;
        _source_stream_matmul_16_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_2230) begin
        _source_stream_matmul_16_source_20_pat_size_3 <= 1;
        _source_stream_matmul_16_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_2230) begin
        _stream_matmul_16_source_20_source_sel <= 3;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_20_source_offset_buf <= _stream_matmul_16_source_20_source_offset;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_count_0 <= _source_stream_matmul_16_source_20_pat_size_0 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_count_1 <= _source_stream_matmul_16_source_20_pat_size_1 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_count_2 <= _source_stream_matmul_16_source_20_pat_size_2 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_count_3 <= _source_stream_matmul_16_source_20_pat_size_3 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_size_buf_0 <= _source_stream_matmul_16_source_20_pat_size_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_size_buf_1 <= _source_stream_matmul_16_source_20_pat_size_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_size_buf_2 <= _source_stream_matmul_16_source_20_pat_size_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_size_buf_3 <= _source_stream_matmul_16_source_20_pat_size_3;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_stride_buf_0 <= _source_stream_matmul_16_source_20_pat_stride_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_stride_buf_1 <= _source_stream_matmul_16_source_20_pat_stride_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_stride_buf_2 <= _source_stream_matmul_16_source_20_pat_stride_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_stride_buf_3 <= _source_stream_matmul_16_source_20_pat_stride_3;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_source_busy && _stream_matmul_16_is_root) begin
        __variable_wdata_2530 <= _stream_matmul_16_source_20_source_ram_rdata;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_20_idle <= 0;
        _stream_matmul_16_source_20_source_ram_raddr <= _stream_matmul_16_source_20_source_pat_all_offset;
        _stream_matmul_16_source_20_source_ram_renable <= 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_0 <= _source_stream_matmul_16_source_20_pat_cur_offset_0 + _source_stream_matmul_16_source_20_pat_stride_buf_0;
        _source_stream_matmul_16_source_20_pat_count_0 <= _source_stream_matmul_16_source_20_pat_count_0 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_16_source_20_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_0 <= 0;
        _source_stream_matmul_16_source_20_pat_count_0 <= _source_stream_matmul_16_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_16_source_20_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_1 <= _source_stream_matmul_16_source_20_pat_cur_offset_1 + _source_stream_matmul_16_source_20_pat_stride_buf_1;
        _source_stream_matmul_16_source_20_pat_count_1 <= _source_stream_matmul_16_source_20_pat_count_1 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_16_source_20_pat_count_0 == 0) && (_source_stream_matmul_16_source_20_pat_count_1 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_1 <= 0;
        _source_stream_matmul_16_source_20_pat_count_1 <= _source_stream_matmul_16_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_16_source_20_pat_count_0 == 0) && (_source_stream_matmul_16_source_20_pat_count_1 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_2 <= _source_stream_matmul_16_source_20_pat_cur_offset_2 + _source_stream_matmul_16_source_20_pat_stride_buf_2;
        _source_stream_matmul_16_source_20_pat_count_2 <= _source_stream_matmul_16_source_20_pat_count_2 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_16_source_20_pat_count_0 == 0) && (_source_stream_matmul_16_source_20_pat_count_1 == 0)) && (_source_stream_matmul_16_source_20_pat_count_2 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_2 <= 0;
        _source_stream_matmul_16_source_20_pat_count_2 <= _source_stream_matmul_16_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_16_source_20_pat_count_0 == 0) && (_source_stream_matmul_16_source_20_pat_count_1 == 0) && (_source_stream_matmul_16_source_20_pat_count_2 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_3 <= _source_stream_matmul_16_source_20_pat_cur_offset_3 + _source_stream_matmul_16_source_20_pat_stride_buf_3;
        _source_stream_matmul_16_source_20_pat_count_3 <= _source_stream_matmul_16_source_20_pat_count_3 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_16_source_20_pat_count_0 == 0) && (_source_stream_matmul_16_source_20_pat_count_1 == 0) && (_source_stream_matmul_16_source_20_pat_count_2 == 0)) && (_source_stream_matmul_16_source_20_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_20_pat_cur_offset_3 <= 0;
        _source_stream_matmul_16_source_20_pat_count_3 <= _source_stream_matmul_16_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 1) && _stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_20_source_ram_renable <= 0;
        _stream_matmul_16_source_20_idle <= 1;
      end 
      if((_stream_matmul_16_source_20_source_pat_fsm_2 == 2) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_20_source_ram_renable <= 0;
        _stream_matmul_16_source_20_idle <= 1;
      end 
      if(_set_flag_2233) begin
        _stream_matmul_16_source_21_source_mode <= 5'b10;
        _stream_matmul_16_source_21_source_offset <= matmul_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_2233) begin
        _source_stream_matmul_16_source_21_pat_size_0 <= cparam_matmul_16_stream_reduce_size;
        _source_stream_matmul_16_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_2233) begin
        _source_stream_matmul_16_source_21_pat_size_1 <= matmul_16_next_stream_num_ops;
        _source_stream_matmul_16_source_21_pat_stride_1 <= cparam_matmul_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_2233) begin
        _source_stream_matmul_16_source_21_pat_size_2 <= 1;
        _source_stream_matmul_16_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_2233) begin
        _source_stream_matmul_16_source_21_pat_size_3 <= 1;
        _source_stream_matmul_16_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_2233) begin
        _stream_matmul_16_source_21_source_sel <= 4;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_21_source_offset_buf <= _stream_matmul_16_source_21_source_offset;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_count_0 <= _source_stream_matmul_16_source_21_pat_size_0 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_count_1 <= _source_stream_matmul_16_source_21_pat_size_1 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_count_2 <= _source_stream_matmul_16_source_21_pat_size_2 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_count_3 <= _source_stream_matmul_16_source_21_pat_size_3 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_size_buf_0 <= _source_stream_matmul_16_source_21_pat_size_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_size_buf_1 <= _source_stream_matmul_16_source_21_pat_size_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_size_buf_2 <= _source_stream_matmul_16_source_21_pat_size_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_size_buf_3 <= _source_stream_matmul_16_source_21_pat_size_3;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_stride_buf_0 <= _source_stream_matmul_16_source_21_pat_stride_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_stride_buf_1 <= _source_stream_matmul_16_source_21_pat_stride_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_stride_buf_2 <= _source_stream_matmul_16_source_21_pat_stride_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_stride_buf_3 <= _source_stream_matmul_16_source_21_pat_stride_3;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_source_busy && _stream_matmul_16_is_root) begin
        __variable_wdata_2551 <= _stream_matmul_16_source_21_source_ram_rdata;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_21_idle <= 0;
        _stream_matmul_16_source_21_source_ram_raddr <= _stream_matmul_16_source_21_source_pat_all_offset;
        _stream_matmul_16_source_21_source_ram_renable <= 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_0 <= _source_stream_matmul_16_source_21_pat_cur_offset_0 + _source_stream_matmul_16_source_21_pat_stride_buf_0;
        _source_stream_matmul_16_source_21_pat_count_0 <= _source_stream_matmul_16_source_21_pat_count_0 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_16_source_21_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_0 <= 0;
        _source_stream_matmul_16_source_21_pat_count_0 <= _source_stream_matmul_16_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_16_source_21_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_1 <= _source_stream_matmul_16_source_21_pat_cur_offset_1 + _source_stream_matmul_16_source_21_pat_stride_buf_1;
        _source_stream_matmul_16_source_21_pat_count_1 <= _source_stream_matmul_16_source_21_pat_count_1 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_16_source_21_pat_count_0 == 0) && (_source_stream_matmul_16_source_21_pat_count_1 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_1 <= 0;
        _source_stream_matmul_16_source_21_pat_count_1 <= _source_stream_matmul_16_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_16_source_21_pat_count_0 == 0) && (_source_stream_matmul_16_source_21_pat_count_1 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_2 <= _source_stream_matmul_16_source_21_pat_cur_offset_2 + _source_stream_matmul_16_source_21_pat_stride_buf_2;
        _source_stream_matmul_16_source_21_pat_count_2 <= _source_stream_matmul_16_source_21_pat_count_2 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_16_source_21_pat_count_0 == 0) && (_source_stream_matmul_16_source_21_pat_count_1 == 0)) && (_source_stream_matmul_16_source_21_pat_count_2 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_2 <= 0;
        _source_stream_matmul_16_source_21_pat_count_2 <= _source_stream_matmul_16_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_16_source_21_pat_count_0 == 0) && (_source_stream_matmul_16_source_21_pat_count_1 == 0) && (_source_stream_matmul_16_source_21_pat_count_2 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_3 <= _source_stream_matmul_16_source_21_pat_cur_offset_3 + _source_stream_matmul_16_source_21_pat_stride_buf_3;
        _source_stream_matmul_16_source_21_pat_count_3 <= _source_stream_matmul_16_source_21_pat_count_3 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_16_source_21_pat_count_0 == 0) && (_source_stream_matmul_16_source_21_pat_count_1 == 0) && (_source_stream_matmul_16_source_21_pat_count_2 == 0)) && (_source_stream_matmul_16_source_21_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_21_pat_cur_offset_3 <= 0;
        _source_stream_matmul_16_source_21_pat_count_3 <= _source_stream_matmul_16_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 1) && _stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_21_source_ram_renable <= 0;
        _stream_matmul_16_source_21_idle <= 1;
      end 
      if((_stream_matmul_16_source_21_source_pat_fsm_3 == 2) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_21_source_ram_renable <= 0;
        _stream_matmul_16_source_21_idle <= 1;
      end 
      if(_set_flag_2236) begin
        _stream_matmul_16_source_22_source_mode <= 5'b10;
        _stream_matmul_16_source_22_source_offset <= matmul_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_2236) begin
        _source_stream_matmul_16_source_22_pat_size_0 <= cparam_matmul_16_stream_reduce_size;
        _source_stream_matmul_16_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_2236) begin
        _source_stream_matmul_16_source_22_pat_size_1 <= matmul_16_next_stream_num_ops;
        _source_stream_matmul_16_source_22_pat_stride_1 <= cparam_matmul_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_2236) begin
        _source_stream_matmul_16_source_22_pat_size_2 <= 1;
        _source_stream_matmul_16_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_2236) begin
        _source_stream_matmul_16_source_22_pat_size_3 <= 1;
        _source_stream_matmul_16_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_2236) begin
        _stream_matmul_16_source_22_source_sel <= 5;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_22_source_offset_buf <= _stream_matmul_16_source_22_source_offset;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_count_0 <= _source_stream_matmul_16_source_22_pat_size_0 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_count_1 <= _source_stream_matmul_16_source_22_pat_size_1 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_count_2 <= _source_stream_matmul_16_source_22_pat_size_2 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_count_3 <= _source_stream_matmul_16_source_22_pat_size_3 - 1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_size_buf_0 <= _source_stream_matmul_16_source_22_pat_size_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_size_buf_1 <= _source_stream_matmul_16_source_22_pat_size_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_size_buf_2 <= _source_stream_matmul_16_source_22_pat_size_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_size_buf_3 <= _source_stream_matmul_16_source_22_pat_size_3;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_stride_buf_0 <= _source_stream_matmul_16_source_22_pat_stride_0;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_stride_buf_1 <= _source_stream_matmul_16_source_22_pat_stride_1;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_stride_buf_2 <= _source_stream_matmul_16_source_22_pat_stride_2;
      end 
      if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_stride_buf_3 <= _source_stream_matmul_16_source_22_pat_stride_3;
      end 
      if(_stream_matmul_16_stream_oready && _stream_matmul_16_source_busy && _stream_matmul_16_is_root) begin
        __variable_wdata_2552 <= _stream_matmul_16_source_22_source_ram_rdata;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_22_idle <= 0;
        _stream_matmul_16_source_22_source_ram_raddr <= _stream_matmul_16_source_22_source_pat_all_offset;
        _stream_matmul_16_source_22_source_ram_renable <= 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_0 <= _source_stream_matmul_16_source_22_pat_cur_offset_0 + _source_stream_matmul_16_source_22_pat_stride_buf_0;
        _source_stream_matmul_16_source_22_pat_count_0 <= _source_stream_matmul_16_source_22_pat_count_0 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && (_source_stream_matmul_16_source_22_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_0 <= 0;
        _source_stream_matmul_16_source_22_pat_count_0 <= _source_stream_matmul_16_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && (_source_stream_matmul_16_source_22_pat_count_0 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_1 <= _source_stream_matmul_16_source_22_pat_cur_offset_1 + _source_stream_matmul_16_source_22_pat_stride_buf_1;
        _source_stream_matmul_16_source_22_pat_count_1 <= _source_stream_matmul_16_source_22_pat_count_1 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && (_source_stream_matmul_16_source_22_pat_count_0 == 0) && (_source_stream_matmul_16_source_22_pat_count_1 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_1 <= 0;
        _source_stream_matmul_16_source_22_pat_count_1 <= _source_stream_matmul_16_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_16_source_22_pat_count_0 == 0) && (_source_stream_matmul_16_source_22_pat_count_1 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_2 <= _source_stream_matmul_16_source_22_pat_cur_offset_2 + _source_stream_matmul_16_source_22_pat_stride_buf_2;
        _source_stream_matmul_16_source_22_pat_count_2 <= _source_stream_matmul_16_source_22_pat_count_2 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_16_source_22_pat_count_0 == 0) && (_source_stream_matmul_16_source_22_pat_count_1 == 0)) && (_source_stream_matmul_16_source_22_pat_count_2 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_2 <= 0;
        _source_stream_matmul_16_source_22_pat_count_2 <= _source_stream_matmul_16_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_16_source_22_pat_count_0 == 0) && (_source_stream_matmul_16_source_22_pat_count_1 == 0) && (_source_stream_matmul_16_source_22_pat_count_2 == 0)) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_3 <= _source_stream_matmul_16_source_22_pat_cur_offset_3 + _source_stream_matmul_16_source_22_pat_stride_buf_3;
        _source_stream_matmul_16_source_22_pat_count_3 <= _source_stream_matmul_16_source_22_pat_count_3 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && ((_source_stream_matmul_16_source_22_pat_count_0 == 0) && (_source_stream_matmul_16_source_22_pat_count_1 == 0) && (_source_stream_matmul_16_source_22_pat_count_2 == 0)) && (_source_stream_matmul_16_source_22_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
        _source_stream_matmul_16_source_22_pat_cur_offset_3 <= 0;
        _source_stream_matmul_16_source_22_pat_count_3 <= _source_stream_matmul_16_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 1) && _stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_22_source_ram_renable <= 0;
        _stream_matmul_16_source_22_idle <= 1;
      end 
      if((_stream_matmul_16_source_22_source_pat_fsm_4 == 2) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_source_22_source_ram_renable <= 0;
        _stream_matmul_16_source_22_idle <= 1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2240 <= _set_flag_2239;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2241 <= _tmp_2240;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2242 <= _tmp_2241;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2243 <= _tmp_2242;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2244 <= _tmp_2243;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2245 <= _tmp_2244;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2246 <= _tmp_2245;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2247 <= _tmp_2246;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2248 <= _tmp_2247;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2249 <= _tmp_2248;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2250 <= _tmp_2249;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2251 <= _tmp_2250;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2252 <= _tmp_2251;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2253 <= _tmp_2252;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2254 <= _tmp_2253;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2255 <= _tmp_2254;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2256 <= _tmp_2255;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2257 <= _tmp_2256;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2258 <= _tmp_2257;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2259 <= _tmp_2258;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2260 <= _tmp_2259;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2261 <= _tmp_2260;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2262 <= _tmp_2261;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2263 <= _tmp_2262;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2264 <= _tmp_2263;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2265 <= _tmp_2264;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2266 <= _tmp_2265;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2267 <= _tmp_2266;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2268 <= _tmp_2267;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2269 <= _tmp_2268;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2270 <= _tmp_2269;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2271 <= _tmp_2270;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2272 <= _tmp_2271;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2273 <= _tmp_2272;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2276 <= _tmp_2275;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2277 <= _tmp_2276;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2278 <= _tmp_2277;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2279 <= _tmp_2278;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2280 <= _tmp_2279;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2281 <= _tmp_2280;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2282 <= _tmp_2281;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2283 <= _tmp_2282;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2284 <= _tmp_2283;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2285 <= _tmp_2284;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2286 <= _tmp_2285;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2287 <= _tmp_2286;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2288 <= _tmp_2287;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2289 <= _tmp_2288;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2290 <= _tmp_2289;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2291 <= _tmp_2290;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2292 <= _tmp_2291;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2293 <= _tmp_2292;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2294 <= _tmp_2293;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2295 <= _tmp_2294;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2296 <= _tmp_2295;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2297 <= _tmp_2296;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2298 <= _tmp_2297;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2299 <= _tmp_2298;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2300 <= _tmp_2299;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2301 <= _tmp_2300;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2302 <= _tmp_2301;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2303 <= _tmp_2302;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2304 <= _tmp_2303;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2305 <= _tmp_2304;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2306 <= _tmp_2305;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2307 <= _tmp_2306;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2308 <= _tmp_2307;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2309 <= _tmp_2308;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2310 <= matmul_16_next_stream_num_ops;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2311 <= _tmp_2310;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2312 <= _tmp_2311;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2313 <= _tmp_2312;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2314 <= _tmp_2313;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2315 <= _tmp_2314;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2316 <= _tmp_2315;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2317 <= _tmp_2316;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2318 <= _tmp_2317;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2319 <= _tmp_2318;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2320 <= _tmp_2319;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2321 <= _tmp_2320;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2322 <= _tmp_2321;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2323 <= _tmp_2322;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2324 <= _tmp_2323;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2325 <= _tmp_2324;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2326 <= _tmp_2325;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2327 <= _tmp_2326;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2328 <= _tmp_2327;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2329 <= _tmp_2328;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2330 <= _tmp_2329;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2331 <= _tmp_2330;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2332 <= _tmp_2331;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2333 <= _tmp_2332;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2334 <= _tmp_2333;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2335 <= _tmp_2334;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2336 <= _tmp_2335;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2337 <= _tmp_2336;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2338 <= _tmp_2337;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2339 <= _tmp_2338;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2340 <= _tmp_2339;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2341 <= _tmp_2340;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2342 <= _tmp_2341;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2343 <= _tmp_2342;
      end 
      if(_tmp_2273) begin
        _stream_matmul_16_sink_33_sink_mode <= 5'b1;
        _stream_matmul_16_sink_33_sink_offset <= _tmp_2309;
        _stream_matmul_16_sink_33_sink_size <= _tmp_2343;
        _stream_matmul_16_sink_33_sink_stride <= 1;
      end 
      if(_tmp_2273) begin
        _stream_matmul_16_sink_33_sink_sel <= 6;
      end 
      if(_stream_matmul_16_sink_start && _stream_matmul_16_sink_33_sink_mode & 5'b1 && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_sink_33_sink_offset_buf <= _stream_matmul_16_sink_33_sink_offset;
        _stream_matmul_16_sink_33_sink_size_buf <= _stream_matmul_16_sink_33_sink_size;
        _stream_matmul_16_sink_33_sink_stride_buf <= _stream_matmul_16_sink_33_sink_stride;
      end 
      if((_stream_matmul_16_sink_33_sink_fsm_5 == 1) && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_sink_33_sink_waddr <= _stream_matmul_16_sink_33_sink_offset_buf - _stream_matmul_16_sink_33_sink_stride_buf;
        _stream_matmul_16_sink_33_sink_count <= _stream_matmul_16_sink_33_sink_size_buf;
      end 
      if((_stream_matmul_16_sink_33_sink_fsm_5 == 2) && stream_matmul_16_sink_34_data && _stream_matmul_16_stream_oready) begin
        _stream_matmul_16_sink_33_sink_waddr <= _stream_matmul_16_sink_33_sink_waddr + _stream_matmul_16_sink_33_sink_stride_buf;
        _stream_matmul_16_sink_33_sink_wdata <= stream_matmul_16_sink_33_data;
        _stream_matmul_16_sink_33_sink_wenable <= 1;
        _stream_matmul_16_sink_33_sink_count <= _stream_matmul_16_sink_33_sink_count - 1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2371 <= _stream_matmul_16_source_start;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2372 <= _tmp_2371;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2373 <= _tmp_2372;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2374 <= _stream_matmul_16_source_start;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2375 <= _tmp_2374;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2376 <= _tmp_2375;
      end 
      if(_stream_matmul_16_stream_oready && _tmp_2376) begin
        __variable_wdata_2450 <= 1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2377 <= _stream_matmul_16_source_start;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2378 <= _tmp_2377;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2379 <= _tmp_2378;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2380 <= _tmp_2379;
      end 
      if(_stream_matmul_16_stream_oready && _tmp_2380) begin
        __variable_wdata_2450 <= 0;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2383 <= _tmp_2382;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2386 <= _tmp_2385;
      end 
      if(_stream_matmul_16_stream_oready && _tmp_2386) begin
        __variable_wdata_2450 <= 1;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2387 <= _stream_matmul_16_source_start;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2388 <= _tmp_2387;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2389 <= _tmp_2388;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2390 <= _tmp_2389;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2391 <= _tmp_2390;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2392 <= _tmp_2391;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2393 <= _tmp_2392;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2394 <= _tmp_2393;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2395 <= _tmp_2394;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2396 <= _tmp_2395;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2397 <= _tmp_2396;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2398 <= _tmp_2397;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2399 <= _tmp_2398;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2400 <= _tmp_2399;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2401 <= _tmp_2400;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2402 <= _tmp_2401;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2403 <= _tmp_2402;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2404 <= _tmp_2403;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2405 <= _tmp_2404;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2406 <= _tmp_2405;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2407 <= _tmp_2406;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2408 <= _tmp_2407;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2409 <= _tmp_2408;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2410 <= _tmp_2409;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2411 <= _tmp_2410;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2412 <= _tmp_2411;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2413 <= _tmp_2412;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2414 <= _tmp_2413;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2415 <= _tmp_2414;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2416 <= _tmp_2415;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2417 <= _tmp_2416;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2418 <= _tmp_2417;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2419 <= _tmp_2418;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2420 <= _tmp_2419;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2421 <= _stream_matmul_16_source_stop;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2422 <= _tmp_2421;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2423 <= _tmp_2422;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2424 <= _tmp_2423;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2425 <= _tmp_2424;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2426 <= _tmp_2425;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2427 <= _tmp_2426;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2428 <= _tmp_2427;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2429 <= _tmp_2428;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2430 <= _tmp_2429;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2431 <= _tmp_2430;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2432 <= _tmp_2431;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2433 <= _tmp_2432;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2434 <= _tmp_2433;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2435 <= _tmp_2434;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2436 <= _tmp_2435;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2437 <= _tmp_2436;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2438 <= _tmp_2437;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2439 <= _tmp_2438;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2440 <= _tmp_2439;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2441 <= _tmp_2440;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2442 <= _tmp_2441;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2443 <= _tmp_2442;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2444 <= _tmp_2443;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2445 <= _tmp_2444;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2446 <= _tmp_2445;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2447 <= _tmp_2446;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2448 <= _tmp_2447;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2449 <= _tmp_2448;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2450 <= _tmp_2449;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2451 <= _tmp_2450;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2452 <= _tmp_2451;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2453 <= _tmp_2452;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2454 <= _tmp_2453;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2455 <= _stream_matmul_16_source_busy;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2456 <= _tmp_2455;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2457 <= _tmp_2456;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2458 <= _tmp_2457;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2459 <= _tmp_2458;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2460 <= _tmp_2459;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2461 <= _tmp_2460;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2462 <= _tmp_2461;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2463 <= _tmp_2462;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2464 <= _tmp_2463;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2465 <= _tmp_2464;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2466 <= _tmp_2465;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2467 <= _tmp_2466;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2468 <= _tmp_2467;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2469 <= _tmp_2468;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2470 <= _tmp_2469;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2471 <= _tmp_2470;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2472 <= _tmp_2471;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2473 <= _tmp_2472;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2474 <= _tmp_2473;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2475 <= _tmp_2474;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2476 <= _tmp_2475;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2477 <= _tmp_2476;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2478 <= _tmp_2477;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2479 <= _tmp_2478;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2480 <= _tmp_2479;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2481 <= _tmp_2480;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2482 <= _tmp_2481;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2483 <= _tmp_2482;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2484 <= _tmp_2483;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2485 <= _tmp_2484;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2486 <= _tmp_2485;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2487 <= _tmp_2486;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2488 <= _tmp_2487;
      end 
      if(_stream_matmul_16_stream_oready) begin
        _tmp_2489 <= _stream_matmul_16_sink_busy;
      end 
      if(!_stream_matmul_16_sink_busy && _tmp_2489) begin
        _stream_matmul_16_busy_reg <= 0;
      end 
      if(_stream_matmul_16_source_busy) begin
        _stream_matmul_16_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_matmul_16_fsm_1 = 1;
  localparam _stream_matmul_16_fsm_2 = 2;
  localparam _stream_matmul_16_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_fsm <= _stream_matmul_16_fsm_init;
      _stream_matmul_16_source_start <= 0;
      _stream_matmul_16_source_busy <= 0;
      _stream_matmul_16_stream_ivalid <= 0;
    end else begin
      if(_stream_matmul_16_stream_oready && _tmp_2373) begin
        _stream_matmul_16_stream_ivalid <= 1;
      end 
      if(_stream_matmul_16_stream_oready && _tmp_2383) begin
        _stream_matmul_16_stream_ivalid <= 0;
      end 
      case(_stream_matmul_16_fsm)
        _stream_matmul_16_fsm_init: begin
          if(_stream_matmul_16_run_flag) begin
            _stream_matmul_16_source_start <= 1;
          end 
          if(_stream_matmul_16_run_flag) begin
            _stream_matmul_16_fsm <= _stream_matmul_16_fsm_1;
          end 
        end
        _stream_matmul_16_fsm_1: begin
          if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_start <= 0;
            _stream_matmul_16_source_busy <= 1;
          end 
          if(_stream_matmul_16_source_start && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_fsm <= _stream_matmul_16_fsm_2;
          end 
        end
        _stream_matmul_16_fsm_2: begin
          if(_stream_matmul_16_stream_oready) begin
            _stream_matmul_16_fsm <= _stream_matmul_16_fsm_3;
          end 
        end
        _stream_matmul_16_fsm_3: begin
          if(_stream_matmul_16_stream_oready && (_stream_matmul_16_source_11_idle && _stream_matmul_16_source_13_idle && _stream_matmul_16_source_15_idle && _stream_matmul_16_source_20_idle && _stream_matmul_16_source_21_idle && _stream_matmul_16_source_22_idle && _stream_matmul_16_source_7_idle && _stream_matmul_16_source_9_idle && (_stream_matmul_16_fsm == 3))) begin
            _stream_matmul_16_source_busy <= 0;
          end 
          if(_stream_matmul_16_stream_oready && (_stream_matmul_16_source_11_idle && _stream_matmul_16_source_13_idle && _stream_matmul_16_source_15_idle && _stream_matmul_16_source_20_idle && _stream_matmul_16_source_21_idle && _stream_matmul_16_source_22_idle && _stream_matmul_16_source_7_idle && _stream_matmul_16_source_9_idle && (_stream_matmul_16_fsm == 3)) && _stream_matmul_16_run_flag) begin
            _stream_matmul_16_source_start <= 1;
          end 
          if(_stream_matmul_16_stream_oready && (_stream_matmul_16_source_11_idle && _stream_matmul_16_source_13_idle && _stream_matmul_16_source_15_idle && _stream_matmul_16_source_20_idle && _stream_matmul_16_source_21_idle && _stream_matmul_16_source_22_idle && _stream_matmul_16_source_7_idle && _stream_matmul_16_source_9_idle && (_stream_matmul_16_fsm == 3))) begin
            _stream_matmul_16_fsm <= _stream_matmul_16_fsm_init;
          end 
          if(_stream_matmul_16_stream_oready && (_stream_matmul_16_source_11_idle && _stream_matmul_16_source_13_idle && _stream_matmul_16_source_15_idle && _stream_matmul_16_source_20_idle && _stream_matmul_16_source_21_idle && _stream_matmul_16_source_22_idle && _stream_matmul_16_source_7_idle && _stream_matmul_16_source_9_idle && (_stream_matmul_16_fsm == 3)) && _stream_matmul_16_run_flag) begin
            _stream_matmul_16_fsm <= _stream_matmul_16_fsm_1;
          end 
        end
      endcase
    end
  end

  localparam main_fsm_1 = 1;
  localparam main_fsm_2 = 2;
  localparam main_fsm_3 = 3;
  localparam main_fsm_4 = 4;
  localparam main_fsm_5 = 5;
  localparam main_fsm_6 = 6;
  localparam main_fsm_7 = 7;
  localparam main_fsm_8 = 8;
  localparam main_fsm_9 = 9;
  localparam main_fsm_10 = 10;
  localparam main_fsm_11 = 11;
  localparam main_fsm_12 = 12;
  localparam main_fsm_13 = 13;
  localparam main_fsm_14 = 14;
  localparam main_fsm_15 = 15;
  localparam main_fsm_16 = 16;
  localparam main_fsm_17 = 17;
  localparam main_fsm_18 = 18;
  localparam main_fsm_19 = 19;
  localparam main_fsm_20 = 20;
  localparam main_fsm_21 = 21;
  localparam main_fsm_22 = 22;
  localparam main_fsm_23 = 23;
  localparam main_fsm_24 = 24;
  localparam main_fsm_25 = 25;
  localparam main_fsm_26 = 26;
  localparam main_fsm_27 = 27;
  localparam main_fsm_28 = 28;
  localparam main_fsm_29 = 29;
  localparam main_fsm_30 = 30;
  localparam main_fsm_31 = 31;
  localparam main_fsm_32 = 32;
  localparam main_fsm_33 = 33;
  localparam main_fsm_34 = 34;
  localparam main_fsm_35 = 35;
  localparam main_fsm_36 = 36;
  localparam main_fsm_37 = 37;
  localparam main_fsm_38 = 38;
  localparam main_fsm_39 = 39;
  localparam main_fsm_40 = 40;
  localparam main_fsm_41 = 41;
  localparam main_fsm_42 = 42;
  localparam main_fsm_43 = 43;
  localparam main_fsm_44 = 44;
  localparam main_fsm_45 = 45;
  localparam main_fsm_46 = 46;
  localparam main_fsm_47 = 47;
  localparam main_fsm_48 = 48;
  localparam main_fsm_49 = 49;
  localparam main_fsm_50 = 50;
  localparam main_fsm_51 = 51;
  localparam main_fsm_52 = 52;
  localparam main_fsm_53 = 53;
  localparam main_fsm_54 = 54;
  localparam main_fsm_55 = 55;
  localparam main_fsm_56 = 56;
  localparam main_fsm_57 = 57;

  always @(posedge CLK) begin
    if(RST) begin
      main_fsm <= main_fsm_init;
      conv2d_4_objaddr <= 0;
      conv2d_4_arg_objaddr_0 <= 0;
      conv2d_4_arg_objaddr_1 <= 0;
      conv2d_4_arg_objaddr_2 <= 0;
      conv2d_4_arg_objaddr_3 <= 0;
      conv2d_4_control_param_index <= 0;
      max_pool_serial_6_objaddr <= 0;
      max_pool_serial_6_arg_objaddr_0 <= 0;
      matmul_16_objaddr <= 0;
      matmul_16_arg_objaddr_0 <= 0;
      matmul_16_arg_objaddr_1 <= 0;
      matmul_16_arg_objaddr_2 <= 0;
      matmul_16_arg_objaddr_3 <= 0;
      matmul_16_control_param_index <= 0;
    end else begin
      case(main_fsm)
        main_fsm_init: begin
          if(_saxi_register_4 != 0) begin
            main_fsm <= main_fsm_1;
          end 
        end
        main_fsm_1: begin
          main_fsm <= main_fsm_2;
        end
        main_fsm_2: begin
          main_fsm <= main_fsm_3;
        end
        main_fsm_3: begin
          main_fsm <= main_fsm_4;
        end
        main_fsm_4: begin
          main_fsm <= main_fsm_5;
        end
        main_fsm_5: begin
          conv2d_4_objaddr <= _saxi_register_33;
          main_fsm <= main_fsm_6;
        end
        main_fsm_6: begin
          conv2d_4_arg_objaddr_0 <= _saxi_register_35;
          main_fsm <= main_fsm_7;
        end
        main_fsm_7: begin
          conv2d_4_arg_objaddr_1 <= _saxi_register_36;
          main_fsm <= main_fsm_8;
        end
        main_fsm_8: begin
          conv2d_4_arg_objaddr_2 <= _saxi_register_36 + 4608;
          main_fsm <= main_fsm_9;
        end
        main_fsm_9: begin
          conv2d_4_arg_objaddr_3 <= _saxi_register_36 + 4736;
          main_fsm <= main_fsm_10;
        end
        main_fsm_10: begin
          conv2d_4_control_param_index <= 0;
          main_fsm <= main_fsm_11;
        end
        main_fsm_11: begin
          main_fsm <= main_fsm_12;
        end
        main_fsm_12: begin
          main_fsm <= main_fsm_13;
        end
        main_fsm_13: begin
          if(control_conv2d_4 == 34) begin
            main_fsm <= main_fsm_14;
          end 
        end
        main_fsm_14: begin
          main_fsm <= main_fsm_15;
        end
        main_fsm_15: begin
          max_pool_serial_6_objaddr <= _saxi_register_33 + 131072;
          main_fsm <= main_fsm_16;
        end
        main_fsm_16: begin
          max_pool_serial_6_arg_objaddr_0 <= _saxi_register_33;
          main_fsm <= main_fsm_17;
        end
        main_fsm_17: begin
          main_fsm <= main_fsm_18;
        end
        main_fsm_18: begin
          main_fsm <= main_fsm_19;
        end
        main_fsm_19: begin
          if(control_max_pool_serial_6 == 19) begin
            main_fsm <= main_fsm_20;
          end 
        end
        main_fsm_20: begin
          main_fsm <= main_fsm_21;
        end
        main_fsm_21: begin
          conv2d_4_objaddr <= _saxi_register_33 + 163840;
          main_fsm <= main_fsm_22;
        end
        main_fsm_22: begin
          conv2d_4_arg_objaddr_0 <= _saxi_register_33 + 131072;
          main_fsm <= main_fsm_23;
        end
        main_fsm_23: begin
          conv2d_4_arg_objaddr_1 <= _saxi_register_36 + 4864;
          main_fsm <= main_fsm_24;
        end
        main_fsm_24: begin
          conv2d_4_arg_objaddr_2 <= _saxi_register_36 + 78592;
          main_fsm <= main_fsm_25;
        end
        main_fsm_25: begin
          conv2d_4_arg_objaddr_3 <= _saxi_register_36 + 78720;
          main_fsm <= main_fsm_26;
        end
        main_fsm_26: begin
          conv2d_4_control_param_index <= 1;
          main_fsm <= main_fsm_27;
        end
        main_fsm_27: begin
          main_fsm <= main_fsm_28;
        end
        main_fsm_28: begin
          main_fsm <= main_fsm_29;
        end
        main_fsm_29: begin
          if(control_conv2d_4 == 34) begin
            main_fsm <= main_fsm_30;
          end 
        end
        main_fsm_30: begin
          main_fsm <= main_fsm_31;
        end
        main_fsm_31: begin
          main_fsm <= main_fsm_32;
        end
        main_fsm_32: begin
          main_fsm <= main_fsm_33;
        end
        main_fsm_33: begin
          matmul_16_objaddr <= _saxi_register_33 + 196608;
          main_fsm <= main_fsm_34;
        end
        main_fsm_34: begin
          matmul_16_arg_objaddr_0 <= _saxi_register_33 + 163840;
          main_fsm <= main_fsm_35;
        end
        main_fsm_35: begin
          matmul_16_arg_objaddr_1 <= _saxi_register_36 + 78848;
          main_fsm <= main_fsm_36;
        end
        main_fsm_36: begin
          matmul_16_arg_objaddr_2 <= _saxi_register_36 + 8467456;
          main_fsm <= main_fsm_37;
        end
        main_fsm_37: begin
          matmul_16_arg_objaddr_3 <= _saxi_register_36 + 8467968;
          main_fsm <= main_fsm_38;
        end
        main_fsm_38: begin
          matmul_16_control_param_index <= 0;
          main_fsm <= main_fsm_39;
        end
        main_fsm_39: begin
          main_fsm <= main_fsm_40;
        end
        main_fsm_40: begin
          main_fsm <= main_fsm_41;
        end
        main_fsm_41: begin
          if(control_matmul_16 == 28) begin
            main_fsm <= main_fsm_42;
          end 
        end
        main_fsm_42: begin
          main_fsm <= main_fsm_43;
        end
        main_fsm_43: begin
          matmul_16_objaddr <= _saxi_register_34;
          main_fsm <= main_fsm_44;
        end
        main_fsm_44: begin
          matmul_16_arg_objaddr_0 <= _saxi_register_33 + 196608;
          main_fsm <= main_fsm_45;
        end
        main_fsm_45: begin
          matmul_16_arg_objaddr_1 <= _saxi_register_36 + 8468480;
          main_fsm <= main_fsm_46;
        end
        main_fsm_46: begin
          matmul_16_arg_objaddr_2 <= _saxi_register_36 + 8473600;
          main_fsm <= main_fsm_47;
        end
        main_fsm_47: begin
          matmul_16_arg_objaddr_3 <= _saxi_register_36 + 8473664;
          main_fsm <= main_fsm_48;
        end
        main_fsm_48: begin
          matmul_16_control_param_index <= 1;
          main_fsm <= main_fsm_49;
        end
        main_fsm_49: begin
          main_fsm <= main_fsm_50;
        end
        main_fsm_50: begin
          main_fsm <= main_fsm_51;
        end
        main_fsm_51: begin
          if(control_matmul_16 == 28) begin
            main_fsm <= main_fsm_52;
          end 
        end
        main_fsm_52: begin
          main_fsm <= main_fsm_53;
        end
        main_fsm_53: begin
          main_fsm <= main_fsm_54;
        end
        main_fsm_54: begin
          main_fsm <= main_fsm_55;
        end
        main_fsm_55: begin
          main_fsm <= main_fsm_56;
        end
        main_fsm_56: begin
          main_fsm <= main_fsm_57;
        end
        main_fsm_57: begin
          main_fsm <= main_fsm_init;
        end
      endcase
    end
  end

  localparam control_conv2d_4_1 = 1;
  localparam control_conv2d_4_2 = 2;
  localparam control_conv2d_4_3 = 3;
  localparam control_conv2d_4_4 = 4;
  localparam control_conv2d_4_5 = 5;
  localparam control_conv2d_4_6 = 6;
  localparam control_conv2d_4_7 = 7;
  localparam control_conv2d_4_8 = 8;
  localparam control_conv2d_4_9 = 9;
  localparam control_conv2d_4_10 = 10;
  localparam control_conv2d_4_11 = 11;
  localparam control_conv2d_4_12 = 12;
  localparam control_conv2d_4_13 = 13;
  localparam control_conv2d_4_14 = 14;
  localparam control_conv2d_4_15 = 15;
  localparam control_conv2d_4_16 = 16;
  localparam control_conv2d_4_17 = 17;
  localparam control_conv2d_4_18 = 18;
  localparam control_conv2d_4_19 = 19;
  localparam control_conv2d_4_20 = 20;
  localparam control_conv2d_4_21 = 21;
  localparam control_conv2d_4_22 = 22;
  localparam control_conv2d_4_23 = 23;
  localparam control_conv2d_4_24 = 24;
  localparam control_conv2d_4_25 = 25;
  localparam control_conv2d_4_26 = 26;
  localparam control_conv2d_4_27 = 27;
  localparam control_conv2d_4_28 = 28;
  localparam control_conv2d_4_29 = 29;
  localparam control_conv2d_4_30 = 30;
  localparam control_conv2d_4_31 = 31;
  localparam control_conv2d_4_32 = 32;
  localparam control_conv2d_4_33 = 33;
  localparam control_conv2d_4_34 = 34;

  always @(posedge CLK) begin
    if(RST) begin
      control_conv2d_4 <= control_conv2d_4_init;
      _control_conv2d_4_called <= 0;
      conv2d_4_filter_base_offset <= 0;
      conv2d_4_filter_page_comp_offset <= 0;
      conv2d_4_filter_page_dma_offset <= 0;
      conv2d_4_act_base_offset_row <= 0;
      conv2d_4_act_base_offset_bat <= 0;
      conv2d_4_dma_flag_0 <= 0;
      conv2d_4_dma_flag_1 <= 0;
      conv2d_4_dma_flag_2 <= 0;
      conv2d_4_act_page_comp_offset_0 <= 0;
      conv2d_4_act_page_comp_offset_1 <= 0;
      conv2d_4_act_page_comp_offset_2 <= 0;
      conv2d_4_act_page_dma_offset_0 <= 0;
      conv2d_4_act_page_dma_offset_1 <= 0;
      conv2d_4_act_page_dma_offset_2 <= 0;
      conv2d_4_out_base_offset_val <= 0;
      conv2d_4_out_base_offset_col <= 0;
      conv2d_4_out_base_offset_row <= 0;
      conv2d_4_out_base_offset_bat <= 0;
      conv2d_4_out_base_offset_och <= 0;
      conv2d_4_out_page <= 0;
      conv2d_4_out_page_comp_offset <= 0;
      conv2d_4_out_page_dma_offset <= 0;
      conv2d_4_out_laddr_offset <= 0;
      conv2d_4_sync_out_count <= 0;
      conv2d_4_write_count <= 0;
      conv2d_4_next_out_write_size <= 0;
      conv2d_4_row_count <= 0;
      conv2d_4_bat_count <= 0;
      conv2d_4_och_count <= 0;
      conv2d_4_row_select <= 0;
      conv2d_4_prev_row_count <= 0;
      conv2d_4_prev_bat_count <= 0;
      conv2d_4_prev_och_count <= 0;
      conv2d_4_prev_row_select <= 0;
      conv2d_4_out_col_count <= 0;
      conv2d_4_out_row_count <= 0;
      conv2d_4_out_ram_select <= 0;
      conv2d_4_skip_read_filter <= 0;
      conv2d_4_skip_read_act <= 0;
      conv2d_4_skip_comp <= 0;
      conv2d_4_skip_write_out <= 1;
    end else begin
      case(control_conv2d_4)
        control_conv2d_4_init: begin
          if(main_fsm == 11) begin
            _control_conv2d_4_called <= 1;
          end 
          if(main_fsm == 27) begin
            _control_conv2d_4_called <= 1;
          end 
          if(main_fsm == 11) begin
            control_conv2d_4 <= control_conv2d_4_1;
          end 
          if(main_fsm == 27) begin
            control_conv2d_4 <= control_conv2d_4_1;
          end 
        end
        control_conv2d_4_1: begin
          control_conv2d_4 <= control_conv2d_4_2;
        end
        control_conv2d_4_2: begin
          conv2d_4_filter_base_offset <= 0;
          conv2d_4_filter_page_comp_offset <= 0;
          conv2d_4_filter_page_dma_offset <= 0;
          conv2d_4_act_base_offset_row <= 0;
          conv2d_4_act_base_offset_bat <= 0;
          conv2d_4_dma_flag_0 <= 1;
          conv2d_4_dma_flag_1 <= 1;
          conv2d_4_dma_flag_2 <= 1;
          conv2d_4_act_page_comp_offset_0 <= 0;
          conv2d_4_act_page_comp_offset_1 <= 0;
          conv2d_4_act_page_comp_offset_2 <= 0;
          conv2d_4_act_page_dma_offset_0 <= 0;
          conv2d_4_act_page_dma_offset_1 <= 0;
          conv2d_4_act_page_dma_offset_2 <= 0;
          conv2d_4_out_base_offset_val <= 0;
          conv2d_4_out_base_offset_col <= 0;
          conv2d_4_out_base_offset_row <= 0;
          conv2d_4_out_base_offset_bat <= 0;
          conv2d_4_out_base_offset_och <= 0;
          conv2d_4_out_page <= 0;
          conv2d_4_out_page_comp_offset <= 0;
          conv2d_4_out_page_dma_offset <= 0;
          conv2d_4_out_laddr_offset <= 0;
          conv2d_4_sync_out_count <= 0;
          conv2d_4_write_count <= 0;
          conv2d_4_next_out_write_size <= (cparam_conv2d_4_max_och_count == 0)? cparam_conv2d_4_out_write_size_res : cparam_conv2d_4_out_write_size;
          conv2d_4_row_count <= 0;
          conv2d_4_bat_count <= 0;
          conv2d_4_och_count <= 0;
          conv2d_4_row_select <= 0;
          conv2d_4_prev_row_count <= 0;
          conv2d_4_prev_bat_count <= 0;
          conv2d_4_prev_och_count <= 0;
          conv2d_4_prev_row_select <= 0;
          conv2d_4_out_col_count <= 0;
          conv2d_4_out_row_count <= 0;
          conv2d_4_out_ram_select <= 0;
          conv2d_4_skip_read_filter <= 0;
          conv2d_4_skip_read_act <= 0;
          conv2d_4_skip_comp <= 0;
          conv2d_4_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_3;
          end 
        end
        control_conv2d_4_3: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_4;
          end 
        end
        control_conv2d_4_4: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_5;
          end 
        end
        control_conv2d_4_5: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_6;
          end 
        end
        control_conv2d_4_6: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
        end
        control_conv2d_4_7: begin
          control_conv2d_4 <= control_conv2d_4_8;
          if(conv2d_4_skip_read_filter) begin
            control_conv2d_4 <= control_conv2d_4_11;
          end 
        end
        control_conv2d_4_8: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_9;
          end 
        end
        control_conv2d_4_9: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_10;
          end 
        end
        control_conv2d_4_10: begin
          control_conv2d_4 <= control_conv2d_4_11;
        end
        control_conv2d_4_11: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_24;
          end 
        end
        control_conv2d_4_12: begin
          control_conv2d_4 <= control_conv2d_4_13;
          if(conv2d_4_skip_read_act) begin
            control_conv2d_4 <= control_conv2d_4_23;
          end 
        end
        control_conv2d_4_13: begin
          control_conv2d_4 <= control_conv2d_4_14;
          if(conv2d_4_mux_dma_pad_mask_0 || !conv2d_4_mux_dma_flag_0) begin
            control_conv2d_4 <= control_conv2d_4_16;
          end 
        end
        control_conv2d_4_14: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_15;
          end 
        end
        control_conv2d_4_15: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_16;
          end 
        end
        control_conv2d_4_16: begin
          control_conv2d_4 <= control_conv2d_4_17;
          if(conv2d_4_mux_dma_pad_mask_1 || !conv2d_4_mux_dma_flag_1) begin
            control_conv2d_4 <= control_conv2d_4_19;
          end 
        end
        control_conv2d_4_17: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_18;
          end 
        end
        control_conv2d_4_18: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_19;
          end 
        end
        control_conv2d_4_19: begin
          control_conv2d_4 <= control_conv2d_4_20;
          if(conv2d_4_mux_dma_pad_mask_2 || !conv2d_4_mux_dma_flag_2) begin
            control_conv2d_4 <= control_conv2d_4_22;
          end 
        end
        control_conv2d_4_20: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_21;
          end 
        end
        control_conv2d_4_21: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_22;
          end 
        end
        control_conv2d_4_22: begin
          control_conv2d_4 <= control_conv2d_4_23;
        end
        control_conv2d_4_23: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_24;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
        end
        control_conv2d_4_24: begin
          if(_maxi_write_idle) begin
            control_conv2d_4 <= control_conv2d_4_25;
          end 
        end
        control_conv2d_4_25: begin
          if(conv2d_4_comp_fsm == 0) begin
            control_conv2d_4 <= control_conv2d_4_26;
          end 
        end
        control_conv2d_4_26: begin
          control_conv2d_4 <= control_conv2d_4_27;
          if(conv2d_4_skip_write_out) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_prev_och_count < cparam_conv2d_4_max_och_count)) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
        end
        control_conv2d_4_27: begin
          if(conv2d_4_sync_comp_count >= conv2d_4_sync_out_count + cparam_conv2d_4_inc_sync_out) begin
            control_conv2d_4 <= control_conv2d_4_28;
          end 
        end
        control_conv2d_4_28: begin
          if(!conv2d_4_dma_out_mask_0) begin
            control_conv2d_4 <= control_conv2d_4_29;
          end 
          if(conv2d_4_dma_out_mask_0) begin
            control_conv2d_4 <= control_conv2d_4_30;
          end 
        end
        control_conv2d_4_29: begin
          if(_maxi_write_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_30;
          end 
        end
        control_conv2d_4_30: begin
          control_conv2d_4 <= control_conv2d_4_31;
        end
        control_conv2d_4_31: begin
          conv2d_4_write_count <= conv2d_4_write_count + 1;
          if(conv2d_4_out_ram_select == 0) begin
            conv2d_4_out_laddr_offset <= conv2d_4_out_laddr_offset + conv2d_4_next_out_write_size;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter) begin
            conv2d_4_out_base_offset_col <= conv2d_4_out_base_offset_col + cparam_conv2d_4_out_col_step;
            conv2d_4_out_col_count <= conv2d_4_out_col_count + 1;
          end 
          conv2d_4_out_ram_select <= conv2d_4_out_ram_select + 1;
          if(conv2d_4_out_ram_select == 0) begin
            conv2d_4_out_ram_select <= 0;
          end 
          conv2d_4_sync_out_count <= conv2d_4_sync_out_count + cparam_conv2d_4_inc_sync_out;
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter && (conv2d_4_write_count >= cparam_conv2d_4_out_num_col - 1) || (cparam_conv2d_4_data_stationary == 0) && cparam_conv2d_4_keep_filter || (cparam_conv2d_4_data_stationary == 1)) begin
            conv2d_4_sync_out_count <= conv2d_4_sync_out_count + (cparam_conv2d_4_inc_sync_out + cparam_conv2d_4_inc_sync_out_res);
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter) begin
            control_conv2d_4 <= control_conv2d_4_26;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter && (conv2d_4_write_count >= cparam_conv2d_4_out_num_col - 1) || (cparam_conv2d_4_data_stationary == 0) && cparam_conv2d_4_keep_filter || (cparam_conv2d_4_data_stationary == 1)) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
        end
        control_conv2d_4_32: begin
          if(conv2d_4_update_filter) begin
            conv2d_4_filter_base_offset <= conv2d_4_filter_base_offset + cparam_conv2d_4_filter_base_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_filter_base_offset <= 0;
          end 
          if(conv2d_4_update_filter) begin
            conv2d_4_och_count <= conv2d_4_och_count + cparam_conv2d_4_och_count_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_och_count <= 0;
          end 
          if(conv2d_4_update_filter) begin
            conv2d_4_filter_page_comp_offset <= conv2d_4_filter_page_comp_offset + cparam_conv2d_4_filter_read_step;
            conv2d_4_filter_page_dma_offset <= conv2d_4_filter_page_dma_offset + cparam_conv2d_4_filter_read_step;
          end 
          if(conv2d_4_update_filter && (conv2d_4_filter_page_comp_offset + cparam_conv2d_4_filter_read_step + cparam_conv2d_4_filter_read_step > 128)) begin
            conv2d_4_filter_page_comp_offset <= 0;
            conv2d_4_filter_page_dma_offset <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_act_base_offset_row <= conv2d_4_act_base_offset_row + cparam_conv2d_4_act_row_step;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_act_base_offset_row <= 0;
            conv2d_4_act_base_offset_bat <= conv2d_4_act_base_offset_bat + cparam_conv2d_4_act_bat_step;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_act_base_offset_bat <= 0;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_0 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_0 <= cparam_conv2d_4_dma_flag_conds_0;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_0 <= 1;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_1 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_1 <= cparam_conv2d_4_dma_flag_conds_1;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_1 <= 1;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_2 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_2 <= cparam_conv2d_4_dma_flag_conds_2;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_2 <= 1;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_row_count <= conv2d_4_row_count + cparam_conv2d_4_stride_row_par_row;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_row_count <= 0;
            conv2d_4_bat_count <= conv2d_4_bat_count + 1;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_bat_count <= 0;
          end 
          if(conv2d_4_update_act && (cparam_conv2d_4_stride_row_par_row < 3)) begin
            conv2d_4_row_select <= conv2d_4_row_select + cparam_conv2d_4_stride_row_par_row;
            conv2d_4_prev_row_select <= conv2d_4_row_select;
          end 
          if(conv2d_4_update_act && (cparam_conv2d_4_stride_row_par_row < 3) && (conv2d_4_row_select + cparam_conv2d_4_stride_row_par_row >= 3)) begin
            conv2d_4_row_select <= conv2d_4_row_select - (3 - cparam_conv2d_4_stride_row_par_row);
            conv2d_4_prev_row_select <= conv2d_4_row_select;
          end 
          if(conv2d_4_update_act && !(cparam_conv2d_4_stride_row_par_row < 3)) begin
            conv2d_4_row_select <= 0;
            conv2d_4_prev_row_select <= 0;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_row_select <= 0;
            conv2d_4_prev_row_select <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_0) begin
            conv2d_4_act_page_comp_offset_0 <= conv2d_4_act_page_comp_offset_0 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_0 <= conv2d_4_act_page_dma_offset_0 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_0 && (conv2d_4_act_page_comp_offset_0 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 512)) begin
            conv2d_4_act_page_comp_offset_0 <= 0;
            conv2d_4_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_0 <= 0;
            conv2d_4_act_page_dma_offset_0 <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_1) begin
            conv2d_4_act_page_comp_offset_1 <= conv2d_4_act_page_comp_offset_1 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_1 <= conv2d_4_act_page_dma_offset_1 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_1 && (conv2d_4_act_page_comp_offset_1 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 512)) begin
            conv2d_4_act_page_comp_offset_1 <= 0;
            conv2d_4_act_page_dma_offset_1 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_1 <= 0;
            conv2d_4_act_page_dma_offset_1 <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_2) begin
            conv2d_4_act_page_comp_offset_2 <= conv2d_4_act_page_comp_offset_2 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_2 <= conv2d_4_act_page_dma_offset_2 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_2 && (conv2d_4_act_page_comp_offset_2 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 512)) begin
            conv2d_4_act_page_comp_offset_2 <= 0;
            conv2d_4_act_page_dma_offset_2 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_2 <= 0;
            conv2d_4_act_page_dma_offset_2 <= 0;
          end 
          conv2d_4_next_out_write_size <= (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)? cparam_conv2d_4_out_write_size_res : cparam_conv2d_4_out_write_size;
          if(!conv2d_4_skip_write_out) begin
            conv2d_4_write_count <= 0;
            conv2d_4_out_laddr_offset <= 0;
            conv2d_4_out_ram_select <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out) begin
            conv2d_4_out_base_offset_col <= 0;
            conv2d_4_out_base_offset_row <= conv2d_4_out_base_offset_row + cparam_conv2d_4_out_row_step;
            conv2d_4_out_col_count <= 0;
            conv2d_4_out_row_count <= conv2d_4_out_row_count + 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_out_base_offset_row <= 0;
            conv2d_4_out_base_offset_bat <= conv2d_4_out_base_offset_bat + cparam_conv2d_4_out_bat_step;
            conv2d_4_out_row_count <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_prev_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_out_base_offset_bat <= 0;
            conv2d_4_out_base_offset_och <= conv2d_4_out_base_offset_och + cparam_conv2d_4_out_och_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_prev_och_count >= cparam_conv2d_4_max_och_count) && !conv2d_4_skip_write_out) begin
            conv2d_4_out_base_offset_row <= conv2d_4_out_base_offset_row + cparam_conv2d_4_out_row_step;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 64;
            conv2d_4_out_page_dma_offset <= 0;
            conv2d_4_out_page <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 0;
            conv2d_4_out_page_dma_offset <= 64;
            conv2d_4_out_page <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) && !conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 64;
            conv2d_4_out_page_dma_offset <= 0;
            conv2d_4_out_page <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) && conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 0;
            conv2d_4_out_page_dma_offset <= 64;
            conv2d_4_out_page <= 0;
          end 
          conv2d_4_prev_row_count <= conv2d_4_row_count;
          conv2d_4_prev_bat_count <= conv2d_4_bat_count;
          conv2d_4_prev_och_count <= conv2d_4_och_count;
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_read_filter <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && cparam_conv2d_4_keep_filter) begin
            conv2d_4_skip_read_filter <= 1;
          end 
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_read_act <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_skip_read_act <= 1;
          end 
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_comp <= 1;
          end 
          if(conv2d_4_skip_write_out && (conv2d_4_prev_row_count == 0) && (conv2d_4_prev_bat_count == 0) && (conv2d_4_prev_och_count == 0)) begin
            conv2d_4_skip_write_out <= 0;
          end 
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if(!conv2d_4_skip_write_out && (conv2d_4_prev_och_count >= cparam_conv2d_4_max_och_count) && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_prev_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            control_conv2d_4 <= control_conv2d_4_33;
          end 
        end
        control_conv2d_4_33: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_conv2d_4 <= control_conv2d_4_34;
          end 
        end
        control_conv2d_4_34: begin
          if(main_fsm == 14) begin
            _control_conv2d_4_called <= 0;
          end 
          if(main_fsm == 30) begin
            _control_conv2d_4_called <= 0;
          end 
          if(main_fsm == 14) begin
            control_conv2d_4 <= control_conv2d_4_init;
          end 
          if(main_fsm == 30) begin
            control_conv2d_4 <= control_conv2d_4_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
      _maxi_read_cont <= 0;
    end else begin
      case(_maxi_read_req_fsm)
        _maxi_read_req_fsm_init: begin
          if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_1;
          end 
        end
        _maxi_read_req_fsm_1: begin
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_cont <= 1;
          end 
          if((maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
            _maxi_read_cont <= 0;
          end 
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_data_fsm_1 = 1;
  localparam _maxi_read_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
    end else begin
      case(_maxi_read_data_fsm)
        _maxi_read_data_fsm_init: begin
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 11)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
        end
        _maxi_read_data_fsm_1: begin
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
        end
        _maxi_read_data_fsm_2: begin
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_0_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_0 <= write_burst_fsm_0_init;
      write_burst_addr_76 <= 0;
      write_burst_stride_77 <= 0;
      write_burst_length_78 <= 0;
      write_burst_done_79 <= 0;
    end else begin
      case(write_burst_fsm_0)
        write_burst_fsm_0_init: begin
          write_burst_addr_76 <= _maxi_read_local_addr_buf;
          write_burst_stride_77 <= _maxi_read_local_stride_buf;
          write_burst_length_78 <= _maxi_read_local_size_buf;
          write_burst_done_79 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_1;
          end 
        end
        write_burst_fsm_0_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_76 <= write_burst_addr_76 + write_burst_stride_77;
            write_burst_length_78 <= write_burst_length_78 - 1;
            write_burst_done_79 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_78 <= 1)) begin
            write_burst_done_79 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_79 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_78 <= 1)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(0) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_1_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_1 <= write_burst_fsm_1_init;
      write_burst_addr_82 <= 0;
      write_burst_stride_83 <= 0;
      write_burst_length_84 <= 0;
      write_burst_done_85 <= 0;
    end else begin
      case(write_burst_fsm_1)
        write_burst_fsm_1_init: begin
          write_burst_addr_82 <= _maxi_read_local_addr_buf;
          write_burst_stride_83 <= _maxi_read_local_stride_buf;
          write_burst_length_84 <= _maxi_read_local_size_buf;
          write_burst_done_85 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_1 <= write_burst_fsm_1_1;
          end 
        end
        write_burst_fsm_1_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_82 <= write_burst_addr_82 + write_burst_stride_83;
            write_burst_length_84 <= write_burst_length_84 - 1;
            write_burst_done_85 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_84 <= 1)) begin
            write_burst_done_85 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_85 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_84 <= 1)) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
          if(0) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_2_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_2 <= write_burst_fsm_2_init;
      write_burst_addr_90 <= 0;
      write_burst_stride_91 <= 0;
      write_burst_length_92 <= 0;
      write_burst_done_93 <= 0;
    end else begin
      case(write_burst_fsm_2)
        write_burst_fsm_2_init: begin
          write_burst_addr_90 <= _maxi_read_local_addr_buf;
          write_burst_stride_91 <= _maxi_read_local_stride_buf;
          write_burst_length_92 <= _maxi_read_local_size_buf;
          write_burst_done_93 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_1;
          end 
        end
        write_burst_fsm_2_1: begin
          if(write_burst_block_ram_wvalid_88) begin
            write_burst_addr_90 <= write_burst_addr_90 + write_burst_stride_91;
            write_burst_length_92 <= write_burst_length_92 - 1;
            write_burst_done_93 <= 0;
          end 
          if(write_burst_block_ram_wvalid_88 && (write_burst_length_92 <= 1)) begin
            write_burst_done_93 <= 1;
          end 
          if(write_burst_block_ram_wvalid_88 && 0) begin
            write_burst_done_93 <= 1;
          end 
          if(write_burst_block_ram_wvalid_88 && (write_burst_length_92 <= 1)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(write_burst_block_ram_wvalid_88 && 0) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(write_burst_block_ram_wquit_89) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_3_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_3 <= write_burst_fsm_3_init;
      write_burst_addr_96 <= 0;
      write_burst_stride_97 <= 0;
      write_burst_length_98 <= 0;
      write_burst_done_99 <= 0;
    end else begin
      case(write_burst_fsm_3)
        write_burst_fsm_3_init: begin
          write_burst_addr_96 <= _maxi_read_local_addr_buf;
          write_burst_stride_97 <= _maxi_read_local_stride_buf;
          write_burst_length_98 <= _maxi_read_local_size_buf;
          write_burst_done_99 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_1;
          end 
        end
        write_burst_fsm_3_1: begin
          if(write_burst_block_ram_wvalid_94) begin
            write_burst_addr_96 <= write_burst_addr_96 + write_burst_stride_97;
            write_burst_length_98 <= write_burst_length_98 - 1;
            write_burst_done_99 <= 0;
          end 
          if(write_burst_block_ram_wvalid_94 && (write_burst_length_98 <= 1)) begin
            write_burst_done_99 <= 1;
          end 
          if(write_burst_block_ram_wvalid_94 && 0) begin
            write_burst_done_99 <= 1;
          end 
          if(write_burst_block_ram_wvalid_94 && (write_burst_length_98 <= 1)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(write_burst_block_ram_wvalid_94 && 0) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(write_burst_block_ram_wquit_95) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_4_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_4 <= write_burst_fsm_4_init;
      write_burst_addr_102 <= 0;
      write_burst_stride_103 <= 0;
      write_burst_length_104 <= 0;
      write_burst_done_105 <= 0;
    end else begin
      case(write_burst_fsm_4)
        write_burst_fsm_4_init: begin
          write_burst_addr_102 <= _maxi_read_local_addr_buf;
          write_burst_stride_103 <= _maxi_read_local_stride_buf;
          write_burst_length_104 <= _maxi_read_local_size_buf;
          write_burst_done_105 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_4 <= write_burst_fsm_4_1;
          end 
        end
        write_burst_fsm_4_1: begin
          if(write_burst_block_ram_wvalid_100) begin
            write_burst_addr_102 <= write_burst_addr_102 + write_burst_stride_103;
            write_burst_length_104 <= write_burst_length_104 - 1;
            write_burst_done_105 <= 0;
          end 
          if(write_burst_block_ram_wvalid_100 && (write_burst_length_104 <= 1)) begin
            write_burst_done_105 <= 1;
          end 
          if(write_burst_block_ram_wvalid_100 && 0) begin
            write_burst_done_105 <= 1;
          end 
          if(write_burst_block_ram_wvalid_100 && (write_burst_length_104 <= 1)) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
          if(write_burst_block_ram_wvalid_100 && 0) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
          if(write_burst_block_ram_wquit_101) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_5_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_5 <= write_burst_fsm_5_init;
      write_burst_addr_108 <= 0;
      write_burst_stride_109 <= 0;
      write_burst_length_110 <= 0;
      write_burst_done_111 <= 0;
    end else begin
      case(write_burst_fsm_5)
        write_burst_fsm_5_init: begin
          write_burst_addr_108 <= _maxi_read_local_addr_buf;
          write_burst_stride_109 <= _maxi_read_local_stride_buf;
          write_burst_length_110 <= _maxi_read_local_size_buf;
          write_burst_done_111 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_5 <= write_burst_fsm_5_1;
          end 
        end
        write_burst_fsm_5_1: begin
          if(write_burst_block_ram_wvalid_106) begin
            write_burst_addr_108 <= write_burst_addr_108 + write_burst_stride_109;
            write_burst_length_110 <= write_burst_length_110 - 1;
            write_burst_done_111 <= 0;
          end 
          if(write_burst_block_ram_wvalid_106 && (write_burst_length_110 <= 1)) begin
            write_burst_done_111 <= 1;
          end 
          if(write_burst_block_ram_wvalid_106 && 0) begin
            write_burst_done_111 <= 1;
          end 
          if(write_burst_block_ram_wvalid_106 && (write_burst_length_110 <= 1)) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
          if(write_burst_block_ram_wvalid_106 && 0) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
          if(write_burst_block_ram_wquit_107) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_6_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_6 <= write_burst_fsm_6_init;
      write_burst_addr_114 <= 0;
      write_burst_stride_115 <= 0;
      write_burst_length_116 <= 0;
      write_burst_done_117 <= 0;
    end else begin
      case(write_burst_fsm_6)
        write_burst_fsm_6_init: begin
          write_burst_addr_114 <= _maxi_read_local_addr_buf;
          write_burst_stride_115 <= _maxi_read_local_stride_buf;
          write_burst_length_116 <= _maxi_read_local_size_buf;
          write_burst_done_117 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_6 <= write_burst_fsm_6_1;
          end 
        end
        write_burst_fsm_6_1: begin
          if(write_burst_block_ram_wvalid_112) begin
            write_burst_addr_114 <= write_burst_addr_114 + write_burst_stride_115;
            write_burst_length_116 <= write_burst_length_116 - 1;
            write_burst_done_117 <= 0;
          end 
          if(write_burst_block_ram_wvalid_112 && (write_burst_length_116 <= 1)) begin
            write_burst_done_117 <= 1;
          end 
          if(write_burst_block_ram_wvalid_112 && 0) begin
            write_burst_done_117 <= 1;
          end 
          if(write_burst_block_ram_wvalid_112 && (write_burst_length_116 <= 1)) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
          if(write_burst_block_ram_wvalid_112 && 0) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
          if(write_burst_block_ram_wquit_113) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_7_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_7 <= write_burst_fsm_7_init;
      write_burst_addr_120 <= 0;
      write_burst_stride_121 <= 0;
      write_burst_length_122 <= 0;
      write_burst_done_123 <= 0;
    end else begin
      case(write_burst_fsm_7)
        write_burst_fsm_7_init: begin
          write_burst_addr_120 <= _maxi_read_local_addr_buf;
          write_burst_stride_121 <= _maxi_read_local_stride_buf;
          write_burst_length_122 <= _maxi_read_local_size_buf;
          write_burst_done_123 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_7 <= write_burst_fsm_7_1;
          end 
        end
        write_burst_fsm_7_1: begin
          if(write_burst_block_ram_wvalid_118) begin
            write_burst_addr_120 <= write_burst_addr_120 + write_burst_stride_121;
            write_burst_length_122 <= write_burst_length_122 - 1;
            write_burst_done_123 <= 0;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_length_122 <= 1)) begin
            write_burst_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_length_122 <= 1)) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
          if(write_burst_block_ram_wquit_119) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_8_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_8 <= write_burst_fsm_8_init;
      write_burst_addr_126 <= 0;
      write_burst_stride_127 <= 0;
      write_burst_length_128 <= 0;
      write_burst_done_129 <= 0;
    end else begin
      case(write_burst_fsm_8)
        write_burst_fsm_8_init: begin
          write_burst_addr_126 <= _maxi_read_local_addr_buf;
          write_burst_stride_127 <= _maxi_read_local_stride_buf;
          write_burst_length_128 <= _maxi_read_local_size_buf;
          write_burst_done_129 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_8 <= write_burst_fsm_8_1;
          end 
        end
        write_burst_fsm_8_1: begin
          if(write_burst_block_ram_wvalid_124) begin
            write_burst_addr_126 <= write_burst_addr_126 + write_burst_stride_127;
            write_burst_length_128 <= write_burst_length_128 - 1;
            write_burst_done_129 <= 0;
          end 
          if(write_burst_block_ram_wvalid_124 && (write_burst_length_128 <= 1)) begin
            write_burst_done_129 <= 1;
          end 
          if(write_burst_block_ram_wvalid_124 && 0) begin
            write_burst_done_129 <= 1;
          end 
          if(write_burst_block_ram_wvalid_124 && (write_burst_length_128 <= 1)) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
          if(write_burst_block_ram_wvalid_124 && 0) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
          if(write_burst_block_ram_wquit_125) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_9_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_9 <= write_burst_fsm_9_init;
      write_burst_addr_132 <= 0;
      write_burst_stride_133 <= 0;
      write_burst_length_134 <= 0;
      write_burst_done_135 <= 0;
    end else begin
      case(write_burst_fsm_9)
        write_burst_fsm_9_init: begin
          write_burst_addr_132 <= _maxi_read_local_addr_buf;
          write_burst_stride_133 <= _maxi_read_local_stride_buf;
          write_burst_length_134 <= _maxi_read_local_size_buf;
          write_burst_done_135 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_9 <= write_burst_fsm_9_1;
          end 
        end
        write_burst_fsm_9_1: begin
          if(write_burst_block_ram_wvalid_130) begin
            write_burst_addr_132 <= write_burst_addr_132 + write_burst_stride_133;
            write_burst_length_134 <= write_burst_length_134 - 1;
            write_burst_done_135 <= 0;
          end 
          if(write_burst_block_ram_wvalid_130 && (write_burst_length_134 <= 1)) begin
            write_burst_done_135 <= 1;
          end 
          if(write_burst_block_ram_wvalid_130 && 0) begin
            write_burst_done_135 <= 1;
          end 
          if(write_burst_block_ram_wvalid_130 && (write_burst_length_134 <= 1)) begin
            write_burst_fsm_9 <= write_burst_fsm_9_init;
          end 
          if(write_burst_block_ram_wvalid_130 && 0) begin
            write_burst_fsm_9 <= write_burst_fsm_9_init;
          end 
          if(write_burst_block_ram_wquit_131) begin
            write_burst_fsm_9 <= write_burst_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_10_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_10 <= write_burst_fsm_10_init;
      write_burst_addr_138 <= 0;
      write_burst_stride_139 <= 0;
      write_burst_length_140 <= 0;
      write_burst_done_141 <= 0;
    end else begin
      case(write_burst_fsm_10)
        write_burst_fsm_10_init: begin
          write_burst_addr_138 <= _maxi_read_local_addr_buf;
          write_burst_stride_139 <= _maxi_read_local_stride_buf;
          write_burst_length_140 <= _maxi_read_local_size_buf;
          write_burst_done_141 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_10 <= write_burst_fsm_10_1;
          end 
        end
        write_burst_fsm_10_1: begin
          if(write_burst_block_ram_wvalid_136) begin
            write_burst_addr_138 <= write_burst_addr_138 + write_burst_stride_139;
            write_burst_length_140 <= write_burst_length_140 - 1;
            write_burst_done_141 <= 0;
          end 
          if(write_burst_block_ram_wvalid_136 && (write_burst_length_140 <= 1)) begin
            write_burst_done_141 <= 1;
          end 
          if(write_burst_block_ram_wvalid_136 && 0) begin
            write_burst_done_141 <= 1;
          end 
          if(write_burst_block_ram_wvalid_136 && (write_burst_length_140 <= 1)) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
          if(write_burst_block_ram_wvalid_136 && 0) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
          if(write_burst_block_ram_wquit_137) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_11_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_11 <= write_burst_fsm_11_init;
      write_burst_addr_144 <= 0;
      write_burst_stride_145 <= 0;
      write_burst_length_146 <= 0;
      write_burst_done_147 <= 0;
    end else begin
      case(write_burst_fsm_11)
        write_burst_fsm_11_init: begin
          write_burst_addr_144 <= _maxi_read_local_addr_buf;
          write_burst_stride_145 <= _maxi_read_local_stride_buf;
          write_burst_length_146 <= _maxi_read_local_size_buf;
          write_burst_done_147 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_11 <= write_burst_fsm_11_1;
          end 
        end
        write_burst_fsm_11_1: begin
          if(write_burst_block_ram_wvalid_142) begin
            write_burst_addr_144 <= write_burst_addr_144 + write_burst_stride_145;
            write_burst_length_146 <= write_burst_length_146 - 1;
            write_burst_done_147 <= 0;
          end 
          if(write_burst_block_ram_wvalid_142 && (write_burst_length_146 <= 1)) begin
            write_burst_done_147 <= 1;
          end 
          if(write_burst_block_ram_wvalid_142 && 0) begin
            write_burst_done_147 <= 1;
          end 
          if(write_burst_block_ram_wvalid_142 && (write_burst_length_146 <= 1)) begin
            write_burst_fsm_11 <= write_burst_fsm_11_init;
          end 
          if(write_burst_block_ram_wvalid_142 && 0) begin
            write_burst_fsm_11 <= write_burst_fsm_11_init;
          end 
          if(write_burst_block_ram_wquit_143) begin
            write_burst_fsm_11 <= write_burst_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_12_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_12 <= write_burst_fsm_12_init;
      write_burst_addr_150 <= 0;
      write_burst_stride_151 <= 0;
      write_burst_length_152 <= 0;
      write_burst_done_153 <= 0;
    end else begin
      case(write_burst_fsm_12)
        write_burst_fsm_12_init: begin
          write_burst_addr_150 <= _maxi_read_local_addr_buf;
          write_burst_stride_151 <= _maxi_read_local_stride_buf;
          write_burst_length_152 <= _maxi_read_local_size_buf;
          write_burst_done_153 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_12 <= write_burst_fsm_12_1;
          end 
        end
        write_burst_fsm_12_1: begin
          if(write_burst_block_ram_wvalid_148) begin
            write_burst_addr_150 <= write_burst_addr_150 + write_burst_stride_151;
            write_burst_length_152 <= write_burst_length_152 - 1;
            write_burst_done_153 <= 0;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_length_152 <= 1)) begin
            write_burst_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_length_152 <= 1)) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
          if(write_burst_block_ram_wquit_149) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_13_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_13 <= write_burst_fsm_13_init;
      write_burst_addr_156 <= 0;
      write_burst_stride_157 <= 0;
      write_burst_length_158 <= 0;
      write_burst_done_159 <= 0;
    end else begin
      case(write_burst_fsm_13)
        write_burst_fsm_13_init: begin
          write_burst_addr_156 <= _maxi_read_local_addr_buf;
          write_burst_stride_157 <= _maxi_read_local_stride_buf;
          write_burst_length_158 <= _maxi_read_local_size_buf;
          write_burst_done_159 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_13 <= write_burst_fsm_13_1;
          end 
        end
        write_burst_fsm_13_1: begin
          if(write_burst_block_ram_wvalid_154) begin
            write_burst_addr_156 <= write_burst_addr_156 + write_burst_stride_157;
            write_burst_length_158 <= write_burst_length_158 - 1;
            write_burst_done_159 <= 0;
          end 
          if(write_burst_block_ram_wvalid_154 && (write_burst_length_158 <= 1)) begin
            write_burst_done_159 <= 1;
          end 
          if(write_burst_block_ram_wvalid_154 && 0) begin
            write_burst_done_159 <= 1;
          end 
          if(write_burst_block_ram_wvalid_154 && (write_burst_length_158 <= 1)) begin
            write_burst_fsm_13 <= write_burst_fsm_13_init;
          end 
          if(write_burst_block_ram_wvalid_154 && 0) begin
            write_burst_fsm_13 <= write_burst_fsm_13_init;
          end 
          if(write_burst_block_ram_wquit_155) begin
            write_burst_fsm_13 <= write_burst_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_14_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_14 <= write_burst_fsm_14_init;
      write_burst_addr_162 <= 0;
      write_burst_stride_163 <= 0;
      write_burst_length_164 <= 0;
      write_burst_done_165 <= 0;
    end else begin
      case(write_burst_fsm_14)
        write_burst_fsm_14_init: begin
          write_burst_addr_162 <= _maxi_read_local_addr_buf;
          write_burst_stride_163 <= _maxi_read_local_stride_buf;
          write_burst_length_164 <= _maxi_read_local_size_buf;
          write_burst_done_165 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_14 <= write_burst_fsm_14_1;
          end 
        end
        write_burst_fsm_14_1: begin
          if(write_burst_block_ram_wvalid_160) begin
            write_burst_addr_162 <= write_burst_addr_162 + write_burst_stride_163;
            write_burst_length_164 <= write_burst_length_164 - 1;
            write_burst_done_165 <= 0;
          end 
          if(write_burst_block_ram_wvalid_160 && (write_burst_length_164 <= 1)) begin
            write_burst_done_165 <= 1;
          end 
          if(write_burst_block_ram_wvalid_160 && 0) begin
            write_burst_done_165 <= 1;
          end 
          if(write_burst_block_ram_wvalid_160 && (write_burst_length_164 <= 1)) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
          if(write_burst_block_ram_wvalid_160 && 0) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
          if(write_burst_block_ram_wquit_161) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_15_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_15 <= write_burst_fsm_15_init;
      write_burst_addr_168 <= 0;
      write_burst_stride_169 <= 0;
      write_burst_length_170 <= 0;
      write_burst_done_171 <= 0;
    end else begin
      case(write_burst_fsm_15)
        write_burst_fsm_15_init: begin
          write_burst_addr_168 <= _maxi_read_local_addr_buf;
          write_burst_stride_169 <= _maxi_read_local_stride_buf;
          write_burst_length_170 <= _maxi_read_local_size_buf;
          write_burst_done_171 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_15 <= write_burst_fsm_15_1;
          end 
        end
        write_burst_fsm_15_1: begin
          if(write_burst_block_ram_wvalid_166) begin
            write_burst_addr_168 <= write_burst_addr_168 + write_burst_stride_169;
            write_burst_length_170 <= write_burst_length_170 - 1;
            write_burst_done_171 <= 0;
          end 
          if(write_burst_block_ram_wvalid_166 && (write_burst_length_170 <= 1)) begin
            write_burst_done_171 <= 1;
          end 
          if(write_burst_block_ram_wvalid_166 && 0) begin
            write_burst_done_171 <= 1;
          end 
          if(write_burst_block_ram_wvalid_166 && (write_burst_length_170 <= 1)) begin
            write_burst_fsm_15 <= write_burst_fsm_15_init;
          end 
          if(write_burst_block_ram_wvalid_166 && 0) begin
            write_burst_fsm_15 <= write_burst_fsm_15_init;
          end 
          if(write_burst_block_ram_wquit_167) begin
            write_burst_fsm_15 <= write_burst_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_16_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_16 <= write_burst_fsm_16_init;
      write_burst_addr_174 <= 0;
      write_burst_stride_175 <= 0;
      write_burst_length_176 <= 0;
      write_burst_done_177 <= 0;
    end else begin
      case(write_burst_fsm_16)
        write_burst_fsm_16_init: begin
          write_burst_addr_174 <= _maxi_read_local_addr_buf;
          write_burst_stride_175 <= _maxi_read_local_stride_buf;
          write_burst_length_176 <= _maxi_read_local_size_buf;
          write_burst_done_177 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_16 <= write_burst_fsm_16_1;
          end 
        end
        write_burst_fsm_16_1: begin
          if(write_burst_block_ram_wvalid_172) begin
            write_burst_addr_174 <= write_burst_addr_174 + write_burst_stride_175;
            write_burst_length_176 <= write_burst_length_176 - 1;
            write_burst_done_177 <= 0;
          end 
          if(write_burst_block_ram_wvalid_172 && (write_burst_length_176 <= 1)) begin
            write_burst_done_177 <= 1;
          end 
          if(write_burst_block_ram_wvalid_172 && 0) begin
            write_burst_done_177 <= 1;
          end 
          if(write_burst_block_ram_wvalid_172 && (write_burst_length_176 <= 1)) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
          if(write_burst_block_ram_wvalid_172 && 0) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
          if(write_burst_block_ram_wquit_173) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_17_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_17 <= write_burst_fsm_17_init;
      write_burst_addr_180 <= 0;
      write_burst_stride_181 <= 0;
      write_burst_length_182 <= 0;
      write_burst_done_183 <= 0;
    end else begin
      case(write_burst_fsm_17)
        write_burst_fsm_17_init: begin
          write_burst_addr_180 <= _maxi_read_local_addr_buf;
          write_burst_stride_181 <= _maxi_read_local_stride_buf;
          write_burst_length_182 <= _maxi_read_local_size_buf;
          write_burst_done_183 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_17 <= write_burst_fsm_17_1;
          end 
        end
        write_burst_fsm_17_1: begin
          if(write_burst_block_ram_wvalid_178) begin
            write_burst_addr_180 <= write_burst_addr_180 + write_burst_stride_181;
            write_burst_length_182 <= write_burst_length_182 - 1;
            write_burst_done_183 <= 0;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_length_182 <= 1)) begin
            write_burst_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_length_182 <= 1)) begin
            write_burst_fsm_17 <= write_burst_fsm_17_init;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_fsm_17 <= write_burst_fsm_17_init;
          end 
          if(write_burst_block_ram_wquit_179) begin
            write_burst_fsm_17 <= write_burst_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_18_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_18 <= write_burst_fsm_18_init;
      write_burst_addr_186 <= 0;
      write_burst_stride_187 <= 0;
      write_burst_length_188 <= 0;
      write_burst_done_189 <= 0;
    end else begin
      case(write_burst_fsm_18)
        write_burst_fsm_18_init: begin
          write_burst_addr_186 <= _maxi_read_local_addr_buf;
          write_burst_stride_187 <= _maxi_read_local_stride_buf;
          write_burst_length_188 <= _maxi_read_local_size_buf;
          write_burst_done_189 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_18 <= write_burst_fsm_18_1;
          end 
        end
        write_burst_fsm_18_1: begin
          if(write_burst_block_ram_wvalid_184) begin
            write_burst_addr_186 <= write_burst_addr_186 + write_burst_stride_187;
            write_burst_length_188 <= write_burst_length_188 - 1;
            write_burst_done_189 <= 0;
          end 
          if(write_burst_block_ram_wvalid_184 && (write_burst_length_188 <= 1)) begin
            write_burst_done_189 <= 1;
          end 
          if(write_burst_block_ram_wvalid_184 && 0) begin
            write_burst_done_189 <= 1;
          end 
          if(write_burst_block_ram_wvalid_184 && (write_burst_length_188 <= 1)) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
          if(write_burst_block_ram_wvalid_184 && 0) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
          if(write_burst_block_ram_wquit_185) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_19_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_19 <= write_burst_fsm_19_init;
      write_burst_addr_192 <= 0;
      write_burst_stride_193 <= 0;
      write_burst_length_194 <= 0;
      write_burst_done_195 <= 0;
    end else begin
      case(write_burst_fsm_19)
        write_burst_fsm_19_init: begin
          write_burst_addr_192 <= _maxi_read_local_addr_buf;
          write_burst_stride_193 <= _maxi_read_local_stride_buf;
          write_burst_length_194 <= _maxi_read_local_size_buf;
          write_burst_done_195 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_19 <= write_burst_fsm_19_1;
          end 
        end
        write_burst_fsm_19_1: begin
          if(write_burst_block_ram_wvalid_190) begin
            write_burst_addr_192 <= write_burst_addr_192 + write_burst_stride_193;
            write_burst_length_194 <= write_burst_length_194 - 1;
            write_burst_done_195 <= 0;
          end 
          if(write_burst_block_ram_wvalid_190 && (write_burst_length_194 <= 1)) begin
            write_burst_done_195 <= 1;
          end 
          if(write_burst_block_ram_wvalid_190 && 0) begin
            write_burst_done_195 <= 1;
          end 
          if(write_burst_block_ram_wvalid_190 && (write_burst_length_194 <= 1)) begin
            write_burst_fsm_19 <= write_burst_fsm_19_init;
          end 
          if(write_burst_block_ram_wvalid_190 && 0) begin
            write_burst_fsm_19 <= write_burst_fsm_19_init;
          end 
          if(write_burst_block_ram_wquit_191) begin
            write_burst_fsm_19 <= write_burst_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_20_1 = 1;
  localparam write_burst_block_fsm_20_2 = 2;
  localparam write_burst_block_fsm_20_3 = 3;
  localparam write_burst_block_fsm_20_4 = 4;
  localparam write_burst_block_fsm_20_5 = 5;
  localparam write_burst_block_fsm_20_6 = 6;
  localparam write_burst_block_fsm_20_7 = 7;
  localparam write_burst_block_fsm_20_8 = 8;
  localparam write_burst_block_fsm_20_9 = 9;
  localparam write_burst_block_fsm_20_10 = 10;
  localparam write_burst_block_fsm_20_11 = 11;
  localparam write_burst_block_fsm_20_12 = 12;
  localparam write_burst_block_fsm_20_13 = 13;
  localparam write_burst_block_fsm_20_14 = 14;
  localparam write_burst_block_fsm_20_15 = 15;
  localparam write_burst_block_fsm_20_16 = 16;
  localparam write_burst_block_fsm_20_17 = 17;
  localparam write_burst_block_fsm_20_18 = 18;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
      write_burst_block_length_196 <= 0;
      write_burst_block_blocksize_197 <= 0;
      write_burst_block_done_198 <= 0;
      write_burst_block_count_199 <= 0;
    end else begin
      case(write_burst_block_fsm_20)
        write_burst_block_fsm_20_init: begin
          write_burst_block_length_196 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_197 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_198 <= 0;
          write_burst_block_count_199 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_1;
          end 
        end
        write_burst_block_fsm_20_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_4;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_4: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_5;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_5: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_6;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_6: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_7;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_7: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_8;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_8: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_9;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_9: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_10;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_10: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_11;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_11: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_12;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_12: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_13;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_13: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_14;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_14: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_15;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_15: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_16;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_16: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_17;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_17: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_18;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
        write_burst_block_fsm_20_18: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_196 <= write_burst_block_length_196 - 1;
            write_burst_block_done_198 <= 0;
            write_burst_block_count_199 <= write_burst_block_count_199 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_198 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_count_199 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_199 == write_burst_block_blocksize_197 - 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_196 <= 1)) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
          if(0) begin
            write_burst_block_fsm_20 <= write_burst_block_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_21_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_21 <= write_burst_fsm_21_init;
      write_burst_addr_204 <= 0;
      write_burst_stride_205 <= 0;
      write_burst_length_206 <= 0;
      write_burst_done_207 <= 0;
    end else begin
      case(write_burst_fsm_21)
        write_burst_fsm_21_init: begin
          write_burst_addr_204 <= _maxi_read_local_addr_buf;
          write_burst_stride_205 <= _maxi_read_local_stride_buf;
          write_burst_length_206 <= _maxi_read_local_size_buf;
          write_burst_done_207 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_21 <= write_burst_fsm_21_1;
          end 
        end
        write_burst_fsm_21_1: begin
          if(write_burst_block_ram_wvalid_202) begin
            write_burst_addr_204 <= write_burst_addr_204 + write_burst_stride_205;
            write_burst_length_206 <= write_burst_length_206 - 1;
            write_burst_done_207 <= 0;
          end 
          if(write_burst_block_ram_wvalid_202 && (write_burst_length_206 <= 1)) begin
            write_burst_done_207 <= 1;
          end 
          if(write_burst_block_ram_wvalid_202 && 0) begin
            write_burst_done_207 <= 1;
          end 
          if(write_burst_block_ram_wvalid_202 && (write_burst_length_206 <= 1)) begin
            write_burst_fsm_21 <= write_burst_fsm_21_init;
          end 
          if(write_burst_block_ram_wvalid_202 && 0) begin
            write_burst_fsm_21 <= write_burst_fsm_21_init;
          end 
          if(write_burst_block_ram_wquit_203) begin
            write_burst_fsm_21 <= write_burst_fsm_21_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_22_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_22 <= write_burst_fsm_22_init;
      write_burst_addr_210 <= 0;
      write_burst_stride_211 <= 0;
      write_burst_length_212 <= 0;
      write_burst_done_213 <= 0;
    end else begin
      case(write_burst_fsm_22)
        write_burst_fsm_22_init: begin
          write_burst_addr_210 <= _maxi_read_local_addr_buf;
          write_burst_stride_211 <= _maxi_read_local_stride_buf;
          write_burst_length_212 <= _maxi_read_local_size_buf;
          write_burst_done_213 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_22 <= write_burst_fsm_22_1;
          end 
        end
        write_burst_fsm_22_1: begin
          if(write_burst_block_ram_wvalid_208) begin
            write_burst_addr_210 <= write_burst_addr_210 + write_burst_stride_211;
            write_burst_length_212 <= write_burst_length_212 - 1;
            write_burst_done_213 <= 0;
          end 
          if(write_burst_block_ram_wvalid_208 && (write_burst_length_212 <= 1)) begin
            write_burst_done_213 <= 1;
          end 
          if(write_burst_block_ram_wvalid_208 && 0) begin
            write_burst_done_213 <= 1;
          end 
          if(write_burst_block_ram_wvalid_208 && (write_burst_length_212 <= 1)) begin
            write_burst_fsm_22 <= write_burst_fsm_22_init;
          end 
          if(write_burst_block_ram_wvalid_208 && 0) begin
            write_burst_fsm_22 <= write_burst_fsm_22_init;
          end 
          if(write_burst_block_ram_wquit_209) begin
            write_burst_fsm_22 <= write_burst_fsm_22_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_23_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_23 <= write_burst_fsm_23_init;
      write_burst_addr_216 <= 0;
      write_burst_stride_217 <= 0;
      write_burst_length_218 <= 0;
      write_burst_done_219 <= 0;
    end else begin
      case(write_burst_fsm_23)
        write_burst_fsm_23_init: begin
          write_burst_addr_216 <= _maxi_read_local_addr_buf;
          write_burst_stride_217 <= _maxi_read_local_stride_buf;
          write_burst_length_218 <= _maxi_read_local_size_buf;
          write_burst_done_219 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_23 <= write_burst_fsm_23_1;
          end 
        end
        write_burst_fsm_23_1: begin
          if(write_burst_block_ram_wvalid_214) begin
            write_burst_addr_216 <= write_burst_addr_216 + write_burst_stride_217;
            write_burst_length_218 <= write_burst_length_218 - 1;
            write_burst_done_219 <= 0;
          end 
          if(write_burst_block_ram_wvalid_214 && (write_burst_length_218 <= 1)) begin
            write_burst_done_219 <= 1;
          end 
          if(write_burst_block_ram_wvalid_214 && 0) begin
            write_burst_done_219 <= 1;
          end 
          if(write_burst_block_ram_wvalid_214 && (write_burst_length_218 <= 1)) begin
            write_burst_fsm_23 <= write_burst_fsm_23_init;
          end 
          if(write_burst_block_ram_wvalid_214 && 0) begin
            write_burst_fsm_23 <= write_burst_fsm_23_init;
          end 
          if(write_burst_block_ram_wquit_215) begin
            write_burst_fsm_23 <= write_burst_fsm_23_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_24_1 = 1;
  localparam write_burst_block_fsm_24_2 = 2;
  localparam write_burst_block_fsm_24_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
      write_burst_block_length_220 <= 0;
      write_burst_block_blocksize_221 <= 0;
      write_burst_block_done_222 <= 0;
      write_burst_block_count_223 <= 0;
    end else begin
      case(write_burst_block_fsm_24)
        write_burst_block_fsm_24_init: begin
          write_burst_block_length_220 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_221 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_222 <= 0;
          write_burst_block_count_223 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_1;
          end 
        end
        write_burst_block_fsm_24_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_220 <= write_burst_block_length_220 - 1;
            write_burst_block_done_222 <= 0;
            write_burst_block_count_223 <= write_burst_block_count_223 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1)) begin
            write_burst_block_done_222 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_222 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_223 == write_burst_block_blocksize_221 - 1)) begin
            write_burst_block_count_223 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_223 == write_burst_block_blocksize_221 - 1)) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1)) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
          if(0) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
        end
        write_burst_block_fsm_24_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_220 <= write_burst_block_length_220 - 1;
            write_burst_block_done_222 <= 0;
            write_burst_block_count_223 <= write_burst_block_count_223 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1)) begin
            write_burst_block_done_222 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_222 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_223 == write_burst_block_blocksize_221 - 1)) begin
            write_burst_block_count_223 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_223 == write_burst_block_blocksize_221 - 1)) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1)) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
          if(0) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
        end
        write_burst_block_fsm_24_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_220 <= write_burst_block_length_220 - 1;
            write_burst_block_done_222 <= 0;
            write_burst_block_count_223 <= write_burst_block_count_223 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1)) begin
            write_burst_block_done_222 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_222 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_223 == write_burst_block_blocksize_221 - 1)) begin
            write_burst_block_count_223 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_223 == write_burst_block_blocksize_221 - 1)) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_220 <= 1)) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
          if(0) begin
            write_burst_block_fsm_24 <= write_burst_block_fsm_24_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_25_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_25 <= write_burst_fsm_25_init;
      write_burst_addr_228 <= 0;
      write_burst_stride_229 <= 0;
      write_burst_length_230 <= 0;
      write_burst_done_231 <= 0;
    end else begin
      case(write_burst_fsm_25)
        write_burst_fsm_25_init: begin
          write_burst_addr_228 <= _maxi_read_local_addr_buf;
          write_burst_stride_229 <= _maxi_read_local_stride_buf;
          write_burst_length_230 <= _maxi_read_local_size_buf;
          write_burst_done_231 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_25 <= write_burst_fsm_25_1;
          end 
        end
        write_burst_fsm_25_1: begin
          if(write_burst_block_ram_wvalid_226) begin
            write_burst_addr_228 <= write_burst_addr_228 + write_burst_stride_229;
            write_burst_length_230 <= write_burst_length_230 - 1;
            write_burst_done_231 <= 0;
          end 
          if(write_burst_block_ram_wvalid_226 && (write_burst_length_230 <= 1)) begin
            write_burst_done_231 <= 1;
          end 
          if(write_burst_block_ram_wvalid_226 && 0) begin
            write_burst_done_231 <= 1;
          end 
          if(write_burst_block_ram_wvalid_226 && (write_burst_length_230 <= 1)) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
          if(write_burst_block_ram_wvalid_226 && 0) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
          if(write_burst_block_ram_wquit_227) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_26_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_26 <= write_burst_fsm_26_init;
      write_burst_addr_234 <= 0;
      write_burst_stride_235 <= 0;
      write_burst_length_236 <= 0;
      write_burst_done_237 <= 0;
    end else begin
      case(write_burst_fsm_26)
        write_burst_fsm_26_init: begin
          write_burst_addr_234 <= _maxi_read_local_addr_buf;
          write_burst_stride_235 <= _maxi_read_local_stride_buf;
          write_burst_length_236 <= _maxi_read_local_size_buf;
          write_burst_done_237 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_26 <= write_burst_fsm_26_1;
          end 
        end
        write_burst_fsm_26_1: begin
          if(write_burst_block_ram_wvalid_232) begin
            write_burst_addr_234 <= write_burst_addr_234 + write_burst_stride_235;
            write_burst_length_236 <= write_burst_length_236 - 1;
            write_burst_done_237 <= 0;
          end 
          if(write_burst_block_ram_wvalid_232 && (write_burst_length_236 <= 1)) begin
            write_burst_done_237 <= 1;
          end 
          if(write_burst_block_ram_wvalid_232 && 0) begin
            write_burst_done_237 <= 1;
          end 
          if(write_burst_block_ram_wvalid_232 && (write_burst_length_236 <= 1)) begin
            write_burst_fsm_26 <= write_burst_fsm_26_init;
          end 
          if(write_burst_block_ram_wvalid_232 && 0) begin
            write_burst_fsm_26 <= write_burst_fsm_26_init;
          end 
          if(write_burst_block_ram_wquit_233) begin
            write_burst_fsm_26 <= write_burst_fsm_26_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_27_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_27 <= write_burst_fsm_27_init;
      write_burst_addr_240 <= 0;
      write_burst_stride_241 <= 0;
      write_burst_length_242 <= 0;
      write_burst_done_243 <= 0;
    end else begin
      case(write_burst_fsm_27)
        write_burst_fsm_27_init: begin
          write_burst_addr_240 <= _maxi_read_local_addr_buf;
          write_burst_stride_241 <= _maxi_read_local_stride_buf;
          write_burst_length_242 <= _maxi_read_local_size_buf;
          write_burst_done_243 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_27 <= write_burst_fsm_27_1;
          end 
        end
        write_burst_fsm_27_1: begin
          if(write_burst_block_ram_wvalid_238) begin
            write_burst_addr_240 <= write_burst_addr_240 + write_burst_stride_241;
            write_burst_length_242 <= write_burst_length_242 - 1;
            write_burst_done_243 <= 0;
          end 
          if(write_burst_block_ram_wvalid_238 && (write_burst_length_242 <= 1)) begin
            write_burst_done_243 <= 1;
          end 
          if(write_burst_block_ram_wvalid_238 && 0) begin
            write_burst_done_243 <= 1;
          end 
          if(write_burst_block_ram_wvalid_238 && (write_burst_length_242 <= 1)) begin
            write_burst_fsm_27 <= write_burst_fsm_27_init;
          end 
          if(write_burst_block_ram_wvalid_238 && 0) begin
            write_burst_fsm_27 <= write_burst_fsm_27_init;
          end 
          if(write_burst_block_ram_wquit_239) begin
            write_burst_fsm_27 <= write_burst_fsm_27_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_28_1 = 1;
  localparam write_burst_block_fsm_28_2 = 2;
  localparam write_burst_block_fsm_28_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
      write_burst_block_length_244 <= 0;
      write_burst_block_blocksize_245 <= 0;
      write_burst_block_done_246 <= 0;
      write_burst_block_count_247 <= 0;
    end else begin
      case(write_burst_block_fsm_28)
        write_burst_block_fsm_28_init: begin
          write_burst_block_length_244 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_245 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_246 <= 0;
          write_burst_block_count_247 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_1;
          end 
        end
        write_burst_block_fsm_28_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_244 <= write_burst_block_length_244 - 1;
            write_burst_block_done_246 <= 0;
            write_burst_block_count_247 <= write_burst_block_count_247 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1)) begin
            write_burst_block_done_246 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_246 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_247 == write_burst_block_blocksize_245 - 1)) begin
            write_burst_block_count_247 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_247 == write_burst_block_blocksize_245 - 1)) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1)) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
          if(0) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
        end
        write_burst_block_fsm_28_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_244 <= write_burst_block_length_244 - 1;
            write_burst_block_done_246 <= 0;
            write_burst_block_count_247 <= write_burst_block_count_247 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1)) begin
            write_burst_block_done_246 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_246 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_247 == write_burst_block_blocksize_245 - 1)) begin
            write_burst_block_count_247 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_247 == write_burst_block_blocksize_245 - 1)) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1)) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
          if(0) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
        end
        write_burst_block_fsm_28_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_244 <= write_burst_block_length_244 - 1;
            write_burst_block_done_246 <= 0;
            write_burst_block_count_247 <= write_burst_block_count_247 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1)) begin
            write_burst_block_done_246 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_246 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_247 == write_burst_block_blocksize_245 - 1)) begin
            write_burst_block_count_247 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_247 == write_burst_block_blocksize_245 - 1)) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_244 <= 1)) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
          if(0) begin
            write_burst_block_fsm_28 <= write_burst_block_fsm_28_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_29_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_29 <= write_burst_fsm_29_init;
      write_burst_addr_252 <= 0;
      write_burst_stride_253 <= 0;
      write_burst_length_254 <= 0;
      write_burst_done_255 <= 0;
    end else begin
      case(write_burst_fsm_29)
        write_burst_fsm_29_init: begin
          write_burst_addr_252 <= _maxi_read_local_addr_buf;
          write_burst_stride_253 <= _maxi_read_local_stride_buf;
          write_burst_length_254 <= _maxi_read_local_size_buf;
          write_burst_done_255 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_29 <= write_burst_fsm_29_1;
          end 
        end
        write_burst_fsm_29_1: begin
          if(write_burst_block_ram_wvalid_250) begin
            write_burst_addr_252 <= write_burst_addr_252 + write_burst_stride_253;
            write_burst_length_254 <= write_burst_length_254 - 1;
            write_burst_done_255 <= 0;
          end 
          if(write_burst_block_ram_wvalid_250 && (write_burst_length_254 <= 1)) begin
            write_burst_done_255 <= 1;
          end 
          if(write_burst_block_ram_wvalid_250 && 0) begin
            write_burst_done_255 <= 1;
          end 
          if(write_burst_block_ram_wvalid_250 && (write_burst_length_254 <= 1)) begin
            write_burst_fsm_29 <= write_burst_fsm_29_init;
          end 
          if(write_burst_block_ram_wvalid_250 && 0) begin
            write_burst_fsm_29 <= write_burst_fsm_29_init;
          end 
          if(write_burst_block_ram_wquit_251) begin
            write_burst_fsm_29 <= write_burst_fsm_29_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_30_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_30 <= write_burst_fsm_30_init;
      write_burst_addr_258 <= 0;
      write_burst_stride_259 <= 0;
      write_burst_length_260 <= 0;
      write_burst_done_261 <= 0;
    end else begin
      case(write_burst_fsm_30)
        write_burst_fsm_30_init: begin
          write_burst_addr_258 <= _maxi_read_local_addr_buf;
          write_burst_stride_259 <= _maxi_read_local_stride_buf;
          write_burst_length_260 <= _maxi_read_local_size_buf;
          write_burst_done_261 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_30 <= write_burst_fsm_30_1;
          end 
        end
        write_burst_fsm_30_1: begin
          if(write_burst_block_ram_wvalid_256) begin
            write_burst_addr_258 <= write_burst_addr_258 + write_burst_stride_259;
            write_burst_length_260 <= write_burst_length_260 - 1;
            write_burst_done_261 <= 0;
          end 
          if(write_burst_block_ram_wvalid_256 && (write_burst_length_260 <= 1)) begin
            write_burst_done_261 <= 1;
          end 
          if(write_burst_block_ram_wvalid_256 && 0) begin
            write_burst_done_261 <= 1;
          end 
          if(write_burst_block_ram_wvalid_256 && (write_burst_length_260 <= 1)) begin
            write_burst_fsm_30 <= write_burst_fsm_30_init;
          end 
          if(write_burst_block_ram_wvalid_256 && 0) begin
            write_burst_fsm_30 <= write_burst_fsm_30_init;
          end 
          if(write_burst_block_ram_wquit_257) begin
            write_burst_fsm_30 <= write_burst_fsm_30_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_31_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_31 <= write_burst_fsm_31_init;
      write_burst_addr_264 <= 0;
      write_burst_stride_265 <= 0;
      write_burst_length_266 <= 0;
      write_burst_done_267 <= 0;
    end else begin
      case(write_burst_fsm_31)
        write_burst_fsm_31_init: begin
          write_burst_addr_264 <= _maxi_read_local_addr_buf;
          write_burst_stride_265 <= _maxi_read_local_stride_buf;
          write_burst_length_266 <= _maxi_read_local_size_buf;
          write_burst_done_267 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_31 <= write_burst_fsm_31_1;
          end 
        end
        write_burst_fsm_31_1: begin
          if(write_burst_block_ram_wvalid_262) begin
            write_burst_addr_264 <= write_burst_addr_264 + write_burst_stride_265;
            write_burst_length_266 <= write_burst_length_266 - 1;
            write_burst_done_267 <= 0;
          end 
          if(write_burst_block_ram_wvalid_262 && (write_burst_length_266 <= 1)) begin
            write_burst_done_267 <= 1;
          end 
          if(write_burst_block_ram_wvalid_262 && 0) begin
            write_burst_done_267 <= 1;
          end 
          if(write_burst_block_ram_wvalid_262 && (write_burst_length_266 <= 1)) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
          if(write_burst_block_ram_wvalid_262 && 0) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
          if(write_burst_block_ram_wquit_263) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_32_1 = 1;
  localparam write_burst_block_fsm_32_2 = 2;
  localparam write_burst_block_fsm_32_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
      write_burst_block_length_268 <= 0;
      write_burst_block_blocksize_269 <= 0;
      write_burst_block_done_270 <= 0;
      write_burst_block_count_271 <= 0;
    end else begin
      case(write_burst_block_fsm_32)
        write_burst_block_fsm_32_init: begin
          write_burst_block_length_268 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_269 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_270 <= 0;
          write_burst_block_count_271 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_1;
          end 
        end
        write_burst_block_fsm_32_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_268 <= write_burst_block_length_268 - 1;
            write_burst_block_done_270 <= 0;
            write_burst_block_count_271 <= write_burst_block_count_271 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1)) begin
            write_burst_block_done_270 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_270 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_271 == write_burst_block_blocksize_269 - 1)) begin
            write_burst_block_count_271 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_271 == write_burst_block_blocksize_269 - 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
        end
        write_burst_block_fsm_32_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_268 <= write_burst_block_length_268 - 1;
            write_burst_block_done_270 <= 0;
            write_burst_block_count_271 <= write_burst_block_count_271 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1)) begin
            write_burst_block_done_270 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_270 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_271 == write_burst_block_blocksize_269 - 1)) begin
            write_burst_block_count_271 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_271 == write_burst_block_blocksize_269 - 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
        end
        write_burst_block_fsm_32_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_268 <= write_burst_block_length_268 - 1;
            write_burst_block_done_270 <= 0;
            write_burst_block_count_271 <= write_burst_block_count_271 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1)) begin
            write_burst_block_done_270 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_270 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_271 == write_burst_block_blocksize_269 - 1)) begin
            write_burst_block_count_271 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_271 == write_burst_block_blocksize_269 - 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_268 <= 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
        end
      endcase
    end
  end

  localparam conv2d_4_comp_fsm_1 = 1;
  localparam conv2d_4_comp_fsm_2 = 2;
  localparam conv2d_4_comp_fsm_3 = 3;
  localparam conv2d_4_comp_fsm_4 = 4;
  localparam conv2d_4_comp_fsm_5 = 5;
  localparam conv2d_4_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      conv2d_4_comp_fsm <= conv2d_4_comp_fsm_init;
      conv2d_4_stream_act_local_0 <= 0;
      conv2d_4_stream_act_local_1 <= 0;
      conv2d_4_stream_act_local_2 <= 0;
      conv2d_4_stream_act_local_3 <= 0;
      conv2d_4_stream_act_local_4 <= 0;
      conv2d_4_stream_act_local_5 <= 0;
      conv2d_4_stream_act_local_6 <= 0;
      conv2d_4_stream_act_local_7 <= 0;
      conv2d_4_stream_act_local_8 <= 0;
      conv2d_4_stream_out_local_col <= 0;
      conv2d_4_stream_out_local_val <= 0;
      conv2d_4_col_count <= 0;
      conv2d_4_col_select <= 0;
      conv2d_4_filter_page_comp_offset_buf <= 0;
      conv2d_4_act_page_comp_offset_buf_0 <= 0;
      conv2d_4_act_page_comp_offset_buf_1 <= 0;
      conv2d_4_act_page_comp_offset_buf_2 <= 0;
      conv2d_4_out_page_comp_offset_buf <= 0;
      conv2d_4_row_count_buf <= 0;
      conv2d_4_row_select_buf <= 0;
      conv2d_4_och_count_buf <= 0;
      conv2d_4_next_stream_num_ops <= 0;
      conv2d_4_stream_pad_masks <= 0;
      conv2d_4_sync_comp_count <= 0;
    end else begin
      if(_stream_conv2d_4_sink_stop) begin
        conv2d_4_sync_comp_count <= conv2d_4_sync_comp_count + 1;
      end 
      if(control_conv2d_4 == 6) begin
        conv2d_4_sync_comp_count <= 0;
      end 
      case(conv2d_4_comp_fsm)
        conv2d_4_comp_fsm_init: begin
          if((control_conv2d_4 == 25) && !conv2d_4_skip_comp) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_1;
          end 
        end
        conv2d_4_comp_fsm_1: begin
          conv2d_4_stream_act_local_0 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_1 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_2 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_3 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_4 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_5 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_6 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_7 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_8 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_out_local_col <= 0;
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count == 0)) begin
            conv2d_4_stream_out_local_val <= 0;
          end 
          conv2d_4_col_count <= 0;
          conv2d_4_col_select <= cparam_conv2d_4_col_select_initval;
          conv2d_4_filter_page_comp_offset_buf <= conv2d_4_filter_page_comp_offset;
          conv2d_4_act_page_comp_offset_buf_0 <= conv2d_4_act_page_comp_offset_0;
          conv2d_4_act_page_comp_offset_buf_1 <= conv2d_4_act_page_comp_offset_1;
          conv2d_4_act_page_comp_offset_buf_2 <= conv2d_4_act_page_comp_offset_2;
          conv2d_4_out_page_comp_offset_buf <= conv2d_4_out_page_comp_offset;
          conv2d_4_row_count_buf <= conv2d_4_row_count;
          conv2d_4_row_select_buf <= conv2d_4_row_select;
          conv2d_4_och_count_buf <= conv2d_4_och_count;
          conv2d_4_next_stream_num_ops <= (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)? cparam_conv2d_4_stream_num_ops_res : cparam_conv2d_4_stream_num_ops;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_2;
        end
        conv2d_4_comp_fsm_2: begin
          conv2d_4_stream_pad_masks <= { conv2d_4_stream_pad_mask_2_2, conv2d_4_stream_pad_mask_2_1, conv2d_4_stream_pad_mask_2_0, conv2d_4_stream_pad_mask_1_2, conv2d_4_stream_pad_mask_1_1, conv2d_4_stream_pad_mask_1_0, conv2d_4_stream_pad_mask_0_2, conv2d_4_stream_pad_mask_0_1, conv2d_4_stream_pad_mask_0_0 };
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_3;
        end
        conv2d_4_comp_fsm_3: begin
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          if(_stream_conv2d_4_stream_oready) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          end 
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
        end
        conv2d_4_comp_fsm_4: begin
          if(!_stream_conv2d_4_source_busy) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_5;
          end 
        end
        conv2d_4_comp_fsm_5: begin
          if(_stream_conv2d_4_busy) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_6;
          end 
        end
        conv2d_4_comp_fsm_6: begin
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_0 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_1 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_2 : 0)) begin
            conv2d_4_stream_act_local_0 <= conv2d_4_stream_act_local_0 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_0 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_1 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_2 : 0) begin
            conv2d_4_stream_act_local_0 <= conv2d_4_stream_act_local_0 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_0 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_3 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_4 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_5 : 0)) begin
            conv2d_4_stream_act_local_1 <= conv2d_4_stream_act_local_1 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_3 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_4 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_5 : 0) begin
            conv2d_4_stream_act_local_1 <= conv2d_4_stream_act_local_1 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_1 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_6 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_7 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_8 : 0)) begin
            conv2d_4_stream_act_local_2 <= conv2d_4_stream_act_local_2 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_6 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_7 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_8 : 0) begin
            conv2d_4_stream_act_local_2 <= conv2d_4_stream_act_local_2 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_2 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_9 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_10 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_11 : 0)) begin
            conv2d_4_stream_act_local_3 <= conv2d_4_stream_act_local_3 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_9 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_10 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_11 : 0) begin
            conv2d_4_stream_act_local_3 <= conv2d_4_stream_act_local_3 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_3 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_12 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_13 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_14 : 0)) begin
            conv2d_4_stream_act_local_4 <= conv2d_4_stream_act_local_4 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_12 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_13 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_14 : 0) begin
            conv2d_4_stream_act_local_4 <= conv2d_4_stream_act_local_4 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_4 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_15 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_16 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_17 : 0)) begin
            conv2d_4_stream_act_local_5 <= conv2d_4_stream_act_local_5 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_15 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_16 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_17 : 0) begin
            conv2d_4_stream_act_local_5 <= conv2d_4_stream_act_local_5 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_5 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_18 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_19 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_20 : 0)) begin
            conv2d_4_stream_act_local_6 <= conv2d_4_stream_act_local_6 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_18 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_19 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_20 : 0) begin
            conv2d_4_stream_act_local_6 <= conv2d_4_stream_act_local_6 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_6 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_21 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_22 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_23 : 0)) begin
            conv2d_4_stream_act_local_7 <= conv2d_4_stream_act_local_7 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_21 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_22 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_23 : 0) begin
            conv2d_4_stream_act_local_7 <= conv2d_4_stream_act_local_7 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_7 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_24 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_25 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_26 : 0)) begin
            conv2d_4_stream_act_local_8 <= conv2d_4_stream_act_local_8 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_24 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_25 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_26 : 0) begin
            conv2d_4_stream_act_local_8 <= conv2d_4_stream_act_local_8 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_8 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(cparam_conv2d_4_data_stationary == 0) begin
            conv2d_4_stream_out_local_col <= conv2d_4_stream_out_local_col + conv2d_4_next_stream_num_ops;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_col_count >= cparam_conv2d_4_max_col_count)) begin
            conv2d_4_stream_out_local_col <= 0;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            conv2d_4_stream_out_local_col <= conv2d_4_stream_out_local_col + cparam_conv2d_4_inc_out_laddr_col;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_col_count >= cparam_conv2d_4_max_col_count)) begin
            conv2d_4_stream_out_local_val <= conv2d_4_stream_out_local_val + conv2d_4_next_stream_num_ops;
            conv2d_4_stream_out_local_col <= 0;
          end 
          conv2d_4_col_count <= conv2d_4_col_count + cparam_conv2d_4_stride_col_par_col;
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_col_count <= 0;
          end 
          conv2d_4_col_select <= conv2d_4_col_select + cparam_conv2d_4_stride_col_mod_filter_num;
          if(conv2d_4_col_select + cparam_conv2d_4_stride_col_mod_filter_num >= 3) begin
            conv2d_4_col_select <= conv2d_4_col_select - cparam_conv2d_4_filter_num_col_minus_stride_col_mod;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_col_select <= cparam_conv2d_4_col_select_initval;
          end 
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_2;
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_conv2d_4_source_7_source_pat_fsm_0)
        _stream_conv2d_4_source_7_source_pat_fsm_0_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_conv2d_4_source_7_source_pat_fsm_0_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0) && (_source_stream_conv2d_4_source_7_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_conv2d_4_source_7_source_pat_fsm_0_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_conv2d_4_source_9_source_pat_fsm_1)
        _stream_conv2d_4_source_9_source_pat_fsm_1_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_conv2d_4_source_9_source_pat_fsm_1_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0) && (_source_stream_conv2d_4_source_9_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_conv2d_4_source_9_source_pat_fsm_1_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_conv2d_4_source_20_source_pat_fsm_2)
        _stream_conv2d_4_source_20_source_pat_fsm_2_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_conv2d_4_source_20_source_pat_fsm_2_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0) && (_source_stream_conv2d_4_source_20_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_conv2d_4_source_20_source_pat_fsm_2_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_conv2d_4_source_21_source_pat_fsm_3)
        _stream_conv2d_4_source_21_source_pat_fsm_3_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_conv2d_4_source_21_source_pat_fsm_3_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0) && (_source_stream_conv2d_4_source_21_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_conv2d_4_source_21_source_pat_fsm_3_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_1 = 1;
  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
    end else begin
      case(_stream_conv2d_4_source_22_source_pat_fsm_4)
        _stream_conv2d_4_source_22_source_pat_fsm_4_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_1;
          end 
        end
        _stream_conv2d_4_source_22_source_pat_fsm_4_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
          end 
          if((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0) && (_source_stream_conv2d_4_source_22_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_2;
          end 
        end
        _stream_conv2d_4_source_22_source_pat_fsm_4_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_1 = 1;
  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
    end else begin
      case(_stream_conv2d_4_source_23_source_pat_fsm_5)
        _stream_conv2d_4_source_23_source_pat_fsm_5_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_1;
          end 
        end
        _stream_conv2d_4_source_23_source_pat_fsm_5_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
          end 
          if((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0) && (_source_stream_conv2d_4_source_23_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_2;
          end 
        end
        _stream_conv2d_4_source_23_source_pat_fsm_5_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_1 = 1;
  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
    end else begin
      case(_stream_conv2d_4_source_24_source_pat_fsm_6)
        _stream_conv2d_4_source_24_source_pat_fsm_6_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_1;
          end 
        end
        _stream_conv2d_4_source_24_source_pat_fsm_6_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
          end 
          if((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0) && (_source_stream_conv2d_4_source_24_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_2;
          end 
        end
        _stream_conv2d_4_source_24_source_pat_fsm_6_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_1 = 1;
  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
    end else begin
      case(_stream_conv2d_4_source_25_source_pat_fsm_7)
        _stream_conv2d_4_source_25_source_pat_fsm_7_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_1;
          end 
        end
        _stream_conv2d_4_source_25_source_pat_fsm_7_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
          end 
          if((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0) && (_source_stream_conv2d_4_source_25_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_2;
          end 
        end
        _stream_conv2d_4_source_25_source_pat_fsm_7_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_1 = 1;
  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
    end else begin
      case(_stream_conv2d_4_source_26_source_pat_fsm_8)
        _stream_conv2d_4_source_26_source_pat_fsm_8_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_1;
          end 
        end
        _stream_conv2d_4_source_26_source_pat_fsm_8_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
          end 
          if((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0) && (_source_stream_conv2d_4_source_26_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_2;
          end 
        end
        _stream_conv2d_4_source_26_source_pat_fsm_8_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_1 = 1;
  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
    end else begin
      case(_stream_conv2d_4_source_27_source_pat_fsm_9)
        _stream_conv2d_4_source_27_source_pat_fsm_9_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_1;
          end 
        end
        _stream_conv2d_4_source_27_source_pat_fsm_9_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
          end 
          if((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0) && (_source_stream_conv2d_4_source_27_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_2;
          end 
        end
        _stream_conv2d_4_source_27_source_pat_fsm_9_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_1 = 1;
  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
    end else begin
      case(_stream_conv2d_4_source_28_source_pat_fsm_10)
        _stream_conv2d_4_source_28_source_pat_fsm_10_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_1;
          end 
        end
        _stream_conv2d_4_source_28_source_pat_fsm_10_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
          end 
          if((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0) && (_source_stream_conv2d_4_source_28_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_2;
          end 
        end
        _stream_conv2d_4_source_28_source_pat_fsm_10_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_1 = 1;
  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
    end else begin
      case(_stream_conv2d_4_source_29_source_pat_fsm_11)
        _stream_conv2d_4_source_29_source_pat_fsm_11_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_1;
          end 
        end
        _stream_conv2d_4_source_29_source_pat_fsm_11_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
          end 
          if((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0) && (_source_stream_conv2d_4_source_29_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_2;
          end 
        end
        _stream_conv2d_4_source_29_source_pat_fsm_11_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_1 = 1;
  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
    end else begin
      case(_stream_conv2d_4_source_30_source_pat_fsm_12)
        _stream_conv2d_4_source_30_source_pat_fsm_12_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_1;
          end 
        end
        _stream_conv2d_4_source_30_source_pat_fsm_12_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
          end 
          if((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0) && (_source_stream_conv2d_4_source_30_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_2;
          end 
        end
        _stream_conv2d_4_source_30_source_pat_fsm_12_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_1 = 1;
  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
    end else begin
      case(_stream_conv2d_4_source_31_source_pat_fsm_13)
        _stream_conv2d_4_source_31_source_pat_fsm_13_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_1;
          end 
        end
        _stream_conv2d_4_source_31_source_pat_fsm_13_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
          end 
          if((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0) && (_source_stream_conv2d_4_source_31_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_2;
          end 
        end
        _stream_conv2d_4_source_31_source_pat_fsm_13_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_1 = 1;
  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
    end else begin
      case(_stream_conv2d_4_source_32_source_pat_fsm_14)
        _stream_conv2d_4_source_32_source_pat_fsm_14_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_1;
          end 
        end
        _stream_conv2d_4_source_32_source_pat_fsm_14_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
          end 
          if((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0) && (_source_stream_conv2d_4_source_32_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_2;
          end 
        end
        _stream_conv2d_4_source_32_source_pat_fsm_14_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_1 = 1;
  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
    end else begin
      case(_stream_conv2d_4_source_33_source_pat_fsm_15)
        _stream_conv2d_4_source_33_source_pat_fsm_15_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_1;
          end 
        end
        _stream_conv2d_4_source_33_source_pat_fsm_15_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
          end 
          if((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0) && (_source_stream_conv2d_4_source_33_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_2;
          end 
        end
        _stream_conv2d_4_source_33_source_pat_fsm_15_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_1 = 1;
  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
    end else begin
      case(_stream_conv2d_4_source_34_source_pat_fsm_16)
        _stream_conv2d_4_source_34_source_pat_fsm_16_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_1;
          end 
        end
        _stream_conv2d_4_source_34_source_pat_fsm_16_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
          end 
          if((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0) && (_source_stream_conv2d_4_source_34_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_2;
          end 
        end
        _stream_conv2d_4_source_34_source_pat_fsm_16_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_1 = 1;
  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
    end else begin
      case(_stream_conv2d_4_source_35_source_pat_fsm_17)
        _stream_conv2d_4_source_35_source_pat_fsm_17_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_1;
          end 
        end
        _stream_conv2d_4_source_35_source_pat_fsm_17_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
          end 
          if((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0) && (_source_stream_conv2d_4_source_35_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_2;
          end 
        end
        _stream_conv2d_4_source_35_source_pat_fsm_17_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_1 = 1;
  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
    end else begin
      case(_stream_conv2d_4_source_36_source_pat_fsm_18)
        _stream_conv2d_4_source_36_source_pat_fsm_18_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_1;
          end 
        end
        _stream_conv2d_4_source_36_source_pat_fsm_18_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
          end 
          if((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0) && (_source_stream_conv2d_4_source_36_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_2;
          end 
        end
        _stream_conv2d_4_source_36_source_pat_fsm_18_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_1 = 1;
  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
    end else begin
      case(_stream_conv2d_4_source_37_source_pat_fsm_19)
        _stream_conv2d_4_source_37_source_pat_fsm_19_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_1;
          end 
        end
        _stream_conv2d_4_source_37_source_pat_fsm_19_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
          end 
          if((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0) && (_source_stream_conv2d_4_source_37_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_2;
          end 
        end
        _stream_conv2d_4_source_37_source_pat_fsm_19_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_38_source_pat_fsm_20_1 = 1;
  localparam _stream_conv2d_4_source_38_source_pat_fsm_20_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_38_source_pat_fsm_20 <= _stream_conv2d_4_source_38_source_pat_fsm_20_init;
    end else begin
      case(_stream_conv2d_4_source_38_source_pat_fsm_20)
        _stream_conv2d_4_source_38_source_pat_fsm_20_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_38_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_38_source_pat_fsm_20 <= _stream_conv2d_4_source_38_source_pat_fsm_20_1;
          end 
        end
        _stream_conv2d_4_source_38_source_pat_fsm_20_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_38_source_pat_fsm_20 <= _stream_conv2d_4_source_38_source_pat_fsm_20_init;
          end 
          if((_source_stream_conv2d_4_source_38_pat_count_0 == 0) && (_source_stream_conv2d_4_source_38_pat_count_1 == 0) && (_source_stream_conv2d_4_source_38_pat_count_2 == 0) && (_source_stream_conv2d_4_source_38_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_38_source_pat_fsm_20 <= _stream_conv2d_4_source_38_source_pat_fsm_20_2;
          end 
        end
        _stream_conv2d_4_source_38_source_pat_fsm_20_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_38_source_pat_fsm_20 <= _stream_conv2d_4_source_38_source_pat_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_39_source_pat_fsm_21_1 = 1;
  localparam _stream_conv2d_4_source_39_source_pat_fsm_21_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_39_source_pat_fsm_21 <= _stream_conv2d_4_source_39_source_pat_fsm_21_init;
    end else begin
      case(_stream_conv2d_4_source_39_source_pat_fsm_21)
        _stream_conv2d_4_source_39_source_pat_fsm_21_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_39_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_39_source_pat_fsm_21 <= _stream_conv2d_4_source_39_source_pat_fsm_21_1;
          end 
        end
        _stream_conv2d_4_source_39_source_pat_fsm_21_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_39_source_pat_fsm_21 <= _stream_conv2d_4_source_39_source_pat_fsm_21_init;
          end 
          if((_source_stream_conv2d_4_source_39_pat_count_0 == 0) && (_source_stream_conv2d_4_source_39_pat_count_1 == 0) && (_source_stream_conv2d_4_source_39_pat_count_2 == 0) && (_source_stream_conv2d_4_source_39_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_39_source_pat_fsm_21 <= _stream_conv2d_4_source_39_source_pat_fsm_21_2;
          end 
        end
        _stream_conv2d_4_source_39_source_pat_fsm_21_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_39_source_pat_fsm_21 <= _stream_conv2d_4_source_39_source_pat_fsm_21_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_40_source_pat_fsm_22_1 = 1;
  localparam _stream_conv2d_4_source_40_source_pat_fsm_22_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_40_source_pat_fsm_22 <= _stream_conv2d_4_source_40_source_pat_fsm_22_init;
    end else begin
      case(_stream_conv2d_4_source_40_source_pat_fsm_22)
        _stream_conv2d_4_source_40_source_pat_fsm_22_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_40_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_40_source_pat_fsm_22 <= _stream_conv2d_4_source_40_source_pat_fsm_22_1;
          end 
        end
        _stream_conv2d_4_source_40_source_pat_fsm_22_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_40_source_pat_fsm_22 <= _stream_conv2d_4_source_40_source_pat_fsm_22_init;
          end 
          if((_source_stream_conv2d_4_source_40_pat_count_0 == 0) && (_source_stream_conv2d_4_source_40_pat_count_1 == 0) && (_source_stream_conv2d_4_source_40_pat_count_2 == 0) && (_source_stream_conv2d_4_source_40_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_40_source_pat_fsm_22 <= _stream_conv2d_4_source_40_source_pat_fsm_22_2;
          end 
        end
        _stream_conv2d_4_source_40_source_pat_fsm_22_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_40_source_pat_fsm_22 <= _stream_conv2d_4_source_40_source_pat_fsm_22_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_41_source_pat_fsm_23_1 = 1;
  localparam _stream_conv2d_4_source_41_source_pat_fsm_23_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_41_source_pat_fsm_23 <= _stream_conv2d_4_source_41_source_pat_fsm_23_init;
    end else begin
      case(_stream_conv2d_4_source_41_source_pat_fsm_23)
        _stream_conv2d_4_source_41_source_pat_fsm_23_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_41_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_41_source_pat_fsm_23 <= _stream_conv2d_4_source_41_source_pat_fsm_23_1;
          end 
        end
        _stream_conv2d_4_source_41_source_pat_fsm_23_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_41_source_pat_fsm_23 <= _stream_conv2d_4_source_41_source_pat_fsm_23_init;
          end 
          if((_source_stream_conv2d_4_source_41_pat_count_0 == 0) && (_source_stream_conv2d_4_source_41_pat_count_1 == 0) && (_source_stream_conv2d_4_source_41_pat_count_2 == 0) && (_source_stream_conv2d_4_source_41_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_41_source_pat_fsm_23 <= _stream_conv2d_4_source_41_source_pat_fsm_23_2;
          end 
        end
        _stream_conv2d_4_source_41_source_pat_fsm_23_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_41_source_pat_fsm_23 <= _stream_conv2d_4_source_41_source_pat_fsm_23_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_42_source_pat_fsm_24_1 = 1;
  localparam _stream_conv2d_4_source_42_source_pat_fsm_24_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_42_source_pat_fsm_24 <= _stream_conv2d_4_source_42_source_pat_fsm_24_init;
    end else begin
      case(_stream_conv2d_4_source_42_source_pat_fsm_24)
        _stream_conv2d_4_source_42_source_pat_fsm_24_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_42_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_42_source_pat_fsm_24 <= _stream_conv2d_4_source_42_source_pat_fsm_24_1;
          end 
        end
        _stream_conv2d_4_source_42_source_pat_fsm_24_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_42_source_pat_fsm_24 <= _stream_conv2d_4_source_42_source_pat_fsm_24_init;
          end 
          if((_source_stream_conv2d_4_source_42_pat_count_0 == 0) && (_source_stream_conv2d_4_source_42_pat_count_1 == 0) && (_source_stream_conv2d_4_source_42_pat_count_2 == 0) && (_source_stream_conv2d_4_source_42_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_42_source_pat_fsm_24 <= _stream_conv2d_4_source_42_source_pat_fsm_24_2;
          end 
        end
        _stream_conv2d_4_source_42_source_pat_fsm_24_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_42_source_pat_fsm_24 <= _stream_conv2d_4_source_42_source_pat_fsm_24_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_43_source_pat_fsm_25_1 = 1;
  localparam _stream_conv2d_4_source_43_source_pat_fsm_25_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_43_source_pat_fsm_25 <= _stream_conv2d_4_source_43_source_pat_fsm_25_init;
    end else begin
      case(_stream_conv2d_4_source_43_source_pat_fsm_25)
        _stream_conv2d_4_source_43_source_pat_fsm_25_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_43_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_43_source_pat_fsm_25 <= _stream_conv2d_4_source_43_source_pat_fsm_25_1;
          end 
        end
        _stream_conv2d_4_source_43_source_pat_fsm_25_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_43_source_pat_fsm_25 <= _stream_conv2d_4_source_43_source_pat_fsm_25_init;
          end 
          if((_source_stream_conv2d_4_source_43_pat_count_0 == 0) && (_source_stream_conv2d_4_source_43_pat_count_1 == 0) && (_source_stream_conv2d_4_source_43_pat_count_2 == 0) && (_source_stream_conv2d_4_source_43_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_43_source_pat_fsm_25 <= _stream_conv2d_4_source_43_source_pat_fsm_25_2;
          end 
        end
        _stream_conv2d_4_source_43_source_pat_fsm_25_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_43_source_pat_fsm_25 <= _stream_conv2d_4_source_43_source_pat_fsm_25_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_44_source_pat_fsm_26_1 = 1;
  localparam _stream_conv2d_4_source_44_source_pat_fsm_26_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_44_source_pat_fsm_26 <= _stream_conv2d_4_source_44_source_pat_fsm_26_init;
    end else begin
      case(_stream_conv2d_4_source_44_source_pat_fsm_26)
        _stream_conv2d_4_source_44_source_pat_fsm_26_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_44_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_44_source_pat_fsm_26 <= _stream_conv2d_4_source_44_source_pat_fsm_26_1;
          end 
        end
        _stream_conv2d_4_source_44_source_pat_fsm_26_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_44_source_pat_fsm_26 <= _stream_conv2d_4_source_44_source_pat_fsm_26_init;
          end 
          if((_source_stream_conv2d_4_source_44_pat_count_0 == 0) && (_source_stream_conv2d_4_source_44_pat_count_1 == 0) && (_source_stream_conv2d_4_source_44_pat_count_2 == 0) && (_source_stream_conv2d_4_source_44_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_44_source_pat_fsm_26 <= _stream_conv2d_4_source_44_source_pat_fsm_26_2;
          end 
        end
        _stream_conv2d_4_source_44_source_pat_fsm_26_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_44_source_pat_fsm_26 <= _stream_conv2d_4_source_44_source_pat_fsm_26_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_45_source_pat_fsm_27_1 = 1;
  localparam _stream_conv2d_4_source_45_source_pat_fsm_27_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_45_source_pat_fsm_27 <= _stream_conv2d_4_source_45_source_pat_fsm_27_init;
    end else begin
      case(_stream_conv2d_4_source_45_source_pat_fsm_27)
        _stream_conv2d_4_source_45_source_pat_fsm_27_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_45_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_45_source_pat_fsm_27 <= _stream_conv2d_4_source_45_source_pat_fsm_27_1;
          end 
        end
        _stream_conv2d_4_source_45_source_pat_fsm_27_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_45_source_pat_fsm_27 <= _stream_conv2d_4_source_45_source_pat_fsm_27_init;
          end 
          if((_source_stream_conv2d_4_source_45_pat_count_0 == 0) && (_source_stream_conv2d_4_source_45_pat_count_1 == 0) && (_source_stream_conv2d_4_source_45_pat_count_2 == 0) && (_source_stream_conv2d_4_source_45_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_45_source_pat_fsm_27 <= _stream_conv2d_4_source_45_source_pat_fsm_27_2;
          end 
        end
        _stream_conv2d_4_source_45_source_pat_fsm_27_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_45_source_pat_fsm_27 <= _stream_conv2d_4_source_45_source_pat_fsm_27_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_source_46_source_pat_fsm_28_1 = 1;
  localparam _stream_conv2d_4_source_46_source_pat_fsm_28_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_46_source_pat_fsm_28 <= _stream_conv2d_4_source_46_source_pat_fsm_28_init;
    end else begin
      case(_stream_conv2d_4_source_46_source_pat_fsm_28)
        _stream_conv2d_4_source_46_source_pat_fsm_28_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_46_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_46_source_pat_fsm_28 <= _stream_conv2d_4_source_46_source_pat_fsm_28_1;
          end 
        end
        _stream_conv2d_4_source_46_source_pat_fsm_28_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_46_source_pat_fsm_28 <= _stream_conv2d_4_source_46_source_pat_fsm_28_init;
          end 
          if((_source_stream_conv2d_4_source_46_pat_count_0 == 0) && (_source_stream_conv2d_4_source_46_pat_count_1 == 0) && (_source_stream_conv2d_4_source_46_pat_count_2 == 0) && (_source_stream_conv2d_4_source_46_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_46_source_pat_fsm_28 <= _stream_conv2d_4_source_46_source_pat_fsm_28_2;
          end 
        end
        _stream_conv2d_4_source_46_source_pat_fsm_28_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_46_source_pat_fsm_28 <= _stream_conv2d_4_source_46_source_pat_fsm_28_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_sink_89_sink_fsm_29_1 = 1;
  localparam _stream_conv2d_4_sink_89_sink_fsm_29_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_sink_89_sink_fsm_29 <= _stream_conv2d_4_sink_89_sink_fsm_29_init;
    end else begin
      case(_stream_conv2d_4_sink_89_sink_fsm_29)
        _stream_conv2d_4_sink_89_sink_fsm_29_init: begin
          if(_stream_conv2d_4_sink_start && _stream_conv2d_4_sink_89_sink_mode & 5'b1 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_89_sink_fsm_29 <= _stream_conv2d_4_sink_89_sink_fsm_29_1;
          end 
        end
        _stream_conv2d_4_sink_89_sink_fsm_29_1: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_89_sink_fsm_29 <= _stream_conv2d_4_sink_89_sink_fsm_29_2;
          end 
        end
        _stream_conv2d_4_sink_89_sink_fsm_29_2: begin
          if(stream_conv2d_4_sink_90_data && (_stream_conv2d_4_sink_89_sink_count == 1) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_89_sink_fsm_29 <= _stream_conv2d_4_sink_89_sink_fsm_29_init;
          end 
          if(_stream_conv2d_4_sink_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_89_sink_fsm_29 <= _stream_conv2d_4_sink_89_sink_fsm_29_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
      _maxi_write_cont <= 0;
    end else begin
      case(_maxi_write_req_fsm)
        _maxi_write_req_fsm_init: begin
          if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_1;
          end 
        end
        _maxi_write_req_fsm_1: begin
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_cont <= 1;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && (_maxi_write_global_size == 0)) begin
            _maxi_write_cont <= 0;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_data_fsm_1 = 1;
  localparam _maxi_write_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
    end else begin
      case(_maxi_write_data_fsm)
        _maxi_write_data_fsm_init: begin
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
        end
        _maxi_write_data_fsm_1: begin
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
        end
        _maxi_write_data_fsm_2: begin
          if((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_2040 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_2041) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_2166 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_2167) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_2495 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_2496) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_33_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_33 <= read_burst_fsm_33_init;
      read_burst_addr_2037 <= 0;
      read_burst_stride_2038 <= 0;
      read_burst_length_2039 <= 0;
      read_burst_rvalid_2040 <= 0;
      read_burst_rlast_2041 <= 0;
    end else begin
      case(read_burst_fsm_33)
        read_burst_fsm_33_init: begin
          read_burst_addr_2037 <= _maxi_write_local_addr_buf;
          read_burst_stride_2038 <= _maxi_write_local_stride_buf;
          read_burst_length_2039 <= _maxi_write_size_buf;
          read_burst_rvalid_2040 <= 0;
          read_burst_rlast_2041 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 1) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_33 <= read_burst_fsm_33_1;
          end 
        end
        read_burst_fsm_33_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2039 > 0)) begin
            read_burst_addr_2037 <= read_burst_addr_2037 + read_burst_stride_2038;
            read_burst_length_2039 <= read_burst_length_2039 - 1;
            read_burst_rvalid_2040 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2039 <= 1)) begin
            read_burst_rlast_2041 <= 1;
          end 
          if(read_burst_rlast_2041 && read_burst_rvalid_2040 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_2040 <= 0;
            read_burst_rlast_2041 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_2040 <= 0;
            read_burst_rlast_2041 <= 0;
          end 
          if(read_burst_rlast_2041 && read_burst_rvalid_2040 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_33 <= read_burst_fsm_33_init;
          end 
          if(0) begin
            read_burst_fsm_33 <= read_burst_fsm_33_init;
          end 
        end
      endcase
    end
  end

  localparam control_max_pool_serial_6_1 = 1;
  localparam control_max_pool_serial_6_2 = 2;
  localparam control_max_pool_serial_6_3 = 3;
  localparam control_max_pool_serial_6_4 = 4;
  localparam control_max_pool_serial_6_5 = 5;
  localparam control_max_pool_serial_6_6 = 6;
  localparam control_max_pool_serial_6_7 = 7;
  localparam control_max_pool_serial_6_8 = 8;
  localparam control_max_pool_serial_6_9 = 9;
  localparam control_max_pool_serial_6_10 = 10;
  localparam control_max_pool_serial_6_11 = 11;
  localparam control_max_pool_serial_6_12 = 12;
  localparam control_max_pool_serial_6_13 = 13;
  localparam control_max_pool_serial_6_14 = 14;
  localparam control_max_pool_serial_6_15 = 15;
  localparam control_max_pool_serial_6_16 = 16;
  localparam control_max_pool_serial_6_17 = 17;
  localparam control_max_pool_serial_6_18 = 18;
  localparam control_max_pool_serial_6_19 = 19;

  always @(posedge CLK) begin
    if(RST) begin
      control_max_pool_serial_6 <= control_max_pool_serial_6_init;
      _control_max_pool_serial_6_called <= 0;
      max_pool_serial_6_act_base_offset_row <= 0;
      max_pool_serial_6_act_base_offset_bat <= 0;
      max_pool_serial_6_act_page <= 0;
      max_pool_serial_6_act_page_comp_offset <= 0;
      max_pool_serial_6_act_page_dma_offset <= 0;
      max_pool_serial_6_out_base_offset_row <= 0;
      max_pool_serial_6_out_base_offset_bat <= 0;
      max_pool_serial_6_out_page <= 0;
      max_pool_serial_6_out_page_comp_offset <= 0;
      max_pool_serial_6_out_page_dma_offset <= 0;
      max_pool_serial_6_row_count <= 0;
      max_pool_serial_6_bat_count <= 0;
      max_pool_serial_6_prev_row_count <= 0;
      max_pool_serial_6_prev_bat_count <= 0;
      max_pool_serial_6_skip_read_act <= 0;
      max_pool_serial_6_skip_comp <= 0;
      max_pool_serial_6_skip_write_out <= 0;
      max_pool_serial_6_out_count <= 0;
    end else begin
      case(control_max_pool_serial_6)
        control_max_pool_serial_6_init: begin
          if(main_fsm == 17) begin
            _control_max_pool_serial_6_called <= 1;
          end 
          if(main_fsm == 17) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_1;
          end 
        end
        control_max_pool_serial_6_1: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_2;
        end
        control_max_pool_serial_6_2: begin
          max_pool_serial_6_act_base_offset_row <= 0;
          max_pool_serial_6_act_base_offset_bat <= 0;
          max_pool_serial_6_act_page <= 0;
          max_pool_serial_6_act_page_comp_offset <= 0;
          max_pool_serial_6_act_page_dma_offset <= 0;
          max_pool_serial_6_out_base_offset_row <= 0;
          max_pool_serial_6_out_base_offset_bat <= 0;
          max_pool_serial_6_out_page <= 0;
          max_pool_serial_6_out_page_comp_offset <= 0;
          max_pool_serial_6_out_page_dma_offset <= 0;
          max_pool_serial_6_row_count <= 0;
          max_pool_serial_6_bat_count <= 0;
          max_pool_serial_6_prev_row_count <= 0;
          max_pool_serial_6_prev_bat_count <= 0;
          max_pool_serial_6_skip_read_act <= 0;
          max_pool_serial_6_skip_comp <= 0;
          max_pool_serial_6_skip_write_out <= 1;
          max_pool_serial_6_out_count <= 0;
          control_max_pool_serial_6 <= control_max_pool_serial_6_3;
        end
        control_max_pool_serial_6_3: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_4;
          if(max_pool_serial_6_skip_read_act) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_11;
          end 
        end
        control_max_pool_serial_6_4: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_5;
          if(max_pool_serial_6_dma_pad_mask_0) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_7;
          end 
        end
        control_max_pool_serial_6_5: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_6;
          end 
        end
        control_max_pool_serial_6_6: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_7;
          end 
        end
        control_max_pool_serial_6_7: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_8;
          if(max_pool_serial_6_dma_pad_mask_1) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_10;
          end 
        end
        control_max_pool_serial_6_8: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_9;
          end 
        end
        control_max_pool_serial_6_9: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_10;
          end 
        end
        control_max_pool_serial_6_10: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_11;
        end
        control_max_pool_serial_6_11: begin
          if(_maxi_write_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_12;
          end 
        end
        control_max_pool_serial_6_12: begin
          if(max_pool_serial_6_comp_fsm == 0) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_13;
          end 
        end
        control_max_pool_serial_6_13: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_14;
          if(max_pool_serial_6_skip_write_out) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_17;
          end 
        end
        control_max_pool_serial_6_14: begin
          if(max_pool_serial_6_comp_count >= max_pool_serial_6_out_count + cparam_max_pool_serial_6_out_write_size) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_15;
          end 
        end
        control_max_pool_serial_6_15: begin
          if(_maxi_write_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_16;
          end 
        end
        control_max_pool_serial_6_16: begin
          max_pool_serial_6_out_count <= max_pool_serial_6_out_count + cparam_max_pool_serial_6_out_write_size;
          control_max_pool_serial_6 <= control_max_pool_serial_6_17;
        end
        control_max_pool_serial_6_17: begin
          max_pool_serial_6_act_base_offset_row <= max_pool_serial_6_act_base_offset_row + cparam_max_pool_serial_6_act_row_step;
          if(max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) begin
            max_pool_serial_6_act_base_offset_row <= 0;
            max_pool_serial_6_act_base_offset_bat <= max_pool_serial_6_act_base_offset_bat + cparam_max_pool_serial_6_act_bat_step;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_act_base_offset_bat <= 0;
          end 
          max_pool_serial_6_row_count <= max_pool_serial_6_row_count + cparam_max_pool_serial_6_stride_row;
          if(max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) begin
            max_pool_serial_6_row_count <= 0;
            max_pool_serial_6_bat_count <= max_pool_serial_6_bat_count + 1;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_bat_count <= 0;
          end 
          if(!max_pool_serial_6_act_page) begin
            max_pool_serial_6_act_page_comp_offset <= 8192;
            max_pool_serial_6_act_page_dma_offset <= 8192;
            max_pool_serial_6_act_page <= 1;
          end 
          if(max_pool_serial_6_act_page) begin
            max_pool_serial_6_act_page_comp_offset <= 0;
            max_pool_serial_6_act_page_dma_offset <= 0;
            max_pool_serial_6_act_page <= 0;
          end 
          if(!max_pool_serial_6_skip_write_out) begin
            max_pool_serial_6_out_base_offset_row <= max_pool_serial_6_out_base_offset_row + cparam_max_pool_serial_6_out_row_step;
          end 
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count)) begin
            max_pool_serial_6_out_base_offset_row <= 0;
            max_pool_serial_6_out_base_offset_bat <= max_pool_serial_6_out_base_offset_bat + cparam_max_pool_serial_6_out_bat_step;
          end 
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_prev_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_out_base_offset_bat <= 0;
          end 
          if(!max_pool_serial_6_out_page) begin
            max_pool_serial_6_out_page_comp_offset <= 4096;
            max_pool_serial_6_out_page_dma_offset <= 0;
            max_pool_serial_6_out_page <= 1;
          end 
          if(max_pool_serial_6_out_page) begin
            max_pool_serial_6_out_page_comp_offset <= 0;
            max_pool_serial_6_out_page_dma_offset <= 4096;
            max_pool_serial_6_out_page <= 0;
          end 
          max_pool_serial_6_prev_row_count <= max_pool_serial_6_row_count;
          max_pool_serial_6_prev_bat_count <= max_pool_serial_6_bat_count;
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_skip_read_act <= 1;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_skip_comp <= 1;
          end 
          if(max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count == 0) && (max_pool_serial_6_prev_bat_count == 0)) begin
            max_pool_serial_6_skip_write_out <= 0;
          end 
          control_max_pool_serial_6 <= control_max_pool_serial_6_3;
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_prev_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_18;
          end 
        end
        control_max_pool_serial_6_18: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_19;
          end 
        end
        control_max_pool_serial_6_19: begin
          if(main_fsm == 20) begin
            _control_max_pool_serial_6_called <= 0;
          end 
          if(main_fsm == 20) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_34_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_34 <= write_burst_fsm_34_init;
      write_burst_addr_2047 <= 0;
      write_burst_stride_2048 <= 0;
      write_burst_length_2049 <= 0;
      write_burst_done_2050 <= 0;
    end else begin
      case(write_burst_fsm_34)
        write_burst_fsm_34_init: begin
          write_burst_addr_2047 <= _maxi_read_local_addr_buf;
          write_burst_stride_2048 <= _maxi_read_local_stride_buf;
          write_burst_length_2049 <= _maxi_read_local_size_buf;
          write_burst_done_2050 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 7) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_34 <= write_burst_fsm_34_1;
          end 
        end
        write_burst_fsm_34_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_2047 <= write_burst_addr_2047 + write_burst_stride_2048;
            write_burst_length_2049 <= write_burst_length_2049 - 1;
            write_burst_done_2050 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2049 <= 1)) begin
            write_burst_done_2050 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_2050 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2049 <= 1)) begin
            write_burst_fsm_34 <= write_burst_fsm_34_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_34 <= write_burst_fsm_34_init;
          end 
          if(0) begin
            write_burst_fsm_34 <= write_burst_fsm_34_init;
          end 
        end
      endcase
    end
  end

  localparam max_pool_serial_6_comp_fsm_1 = 1;
  localparam max_pool_serial_6_comp_fsm_2 = 2;
  localparam max_pool_serial_6_comp_fsm_3 = 3;
  localparam max_pool_serial_6_comp_fsm_4 = 4;
  localparam max_pool_serial_6_comp_fsm_5 = 5;
  localparam max_pool_serial_6_comp_fsm_6 = 6;
  localparam max_pool_serial_6_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_init;
      max_pool_serial_6_stream_act_local <= 0;
      max_pool_serial_6_stream_out_local <= 0;
      max_pool_serial_6_col_count <= 0;
      max_pool_serial_6_act_page_comp_offset_buf <= 0;
      max_pool_serial_6_out_page_comp_offset_buf <= 0;
      max_pool_serial_6_row_count_buf <= 0;
      max_pool_serial_6_stream_pad_masks <= 0;
      max_pool_serial_6_comp_count <= 0;
    end else begin
      if(control_max_pool_serial_6 == 2) begin
        max_pool_serial_6_comp_count <= 0;
      end 
      if(_stream_max_pool_serial_6_sink_stop) begin
        max_pool_serial_6_comp_count <= max_pool_serial_6_comp_count + cparam_max_pool_serial_6_inc_out_laddr;
      end 
      case(max_pool_serial_6_comp_fsm)
        max_pool_serial_6_comp_fsm_init: begin
          if((control_max_pool_serial_6 == 12) && !max_pool_serial_6_skip_comp) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_1;
          end 
        end
        max_pool_serial_6_comp_fsm_1: begin
          max_pool_serial_6_stream_act_local <= cparam_max_pool_serial_6_local_pad_offset;
          max_pool_serial_6_stream_out_local <= 0;
          max_pool_serial_6_col_count <= 0;
          max_pool_serial_6_act_page_comp_offset_buf <= max_pool_serial_6_act_page_comp_offset;
          max_pool_serial_6_out_page_comp_offset_buf <= max_pool_serial_6_out_page_comp_offset;
          max_pool_serial_6_row_count_buf <= max_pool_serial_6_row_count;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_2;
        end
        max_pool_serial_6_comp_fsm_2: begin
          max_pool_serial_6_stream_pad_masks <= { max_pool_serial_6_stream_pad_mask_1_1, max_pool_serial_6_stream_pad_mask_1_0, max_pool_serial_6_stream_pad_mask_0_1, max_pool_serial_6_stream_pad_mask_0_0 };
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_3;
        end
        max_pool_serial_6_comp_fsm_3: begin
          if(!_stream_max_pool_serial_6_source_busy) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_4;
          end 
        end
        max_pool_serial_6_comp_fsm_4: begin
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          if(_stream_max_pool_serial_6_stream_oready) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          end 
        end
        max_pool_serial_6_comp_fsm_5: begin
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_6;
        end
        max_pool_serial_6_comp_fsm_6: begin
          if(_stream_max_pool_serial_6_busy) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_7;
          end 
        end
        max_pool_serial_6_comp_fsm_7: begin
          max_pool_serial_6_stream_act_local <= max_pool_serial_6_stream_act_local + cparam_max_pool_serial_6_inc_act_laddr;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_stream_act_local <= cparam_max_pool_serial_6_local_pad_offset;
          end 
          max_pool_serial_6_stream_out_local <= max_pool_serial_6_stream_out_local + cparam_max_pool_serial_6_inc_out_laddr;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_stream_out_local <= 0;
          end 
          max_pool_serial_6_col_count <= max_pool_serial_6_col_count + cparam_max_pool_serial_6_stride_col;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_col_count <= 0;
          end 
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_2;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1 = 1;
  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
    end else begin
      case(_stream_max_pool_serial_6_source_1_source_pat_fsm_0)
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init: begin
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1;
          end 
        end
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1: begin
          if(_stream_max_pool_serial_6_source_stop && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
          end 
          if((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_3 == 0) && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2;
          end 
        end
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_6_sink_6_sink_fsm_1_1 = 1;
  localparam _stream_max_pool_serial_6_sink_6_sink_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_init;
    end else begin
      case(_stream_max_pool_serial_6_sink_6_sink_fsm_1)
        _stream_max_pool_serial_6_sink_6_sink_fsm_1_init: begin
          if(_stream_max_pool_serial_6_sink_start && _stream_max_pool_serial_6_sink_6_sink_mode & 5'b1 && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_1;
          end 
        end
        _stream_max_pool_serial_6_sink_6_sink_fsm_1_1: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_2;
          end 
        end
        _stream_max_pool_serial_6_sink_6_sink_fsm_1_2: begin
          if(stream_max_pool_serial_6_sink_7_data && (_stream_max_pool_serial_6_sink_6_sink_count == 1) && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_init;
          end 
          if(_stream_max_pool_serial_6_sink_stop && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_6_sink_fsm_1 <= _stream_max_pool_serial_6_sink_6_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_35_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_35 <= read_burst_fsm_35_init;
      read_burst_addr_2163 <= 0;
      read_burst_stride_2164 <= 0;
      read_burst_length_2165 <= 0;
      read_burst_rvalid_2166 <= 0;
      read_burst_rlast_2167 <= 0;
    end else begin
      case(read_burst_fsm_35)
        read_burst_fsm_35_init: begin
          read_burst_addr_2163 <= _maxi_write_local_addr_buf;
          read_burst_stride_2164 <= _maxi_write_local_stride_buf;
          read_burst_length_2165 <= _maxi_write_size_buf;
          read_burst_rvalid_2166 <= 0;
          read_burst_rlast_2167 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 2) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_35 <= read_burst_fsm_35_1;
          end 
        end
        read_burst_fsm_35_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2165 > 0)) begin
            read_burst_addr_2163 <= read_burst_addr_2163 + read_burst_stride_2164;
            read_burst_length_2165 <= read_burst_length_2165 - 1;
            read_burst_rvalid_2166 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2165 <= 1)) begin
            read_burst_rlast_2167 <= 1;
          end 
          if(read_burst_rlast_2167 && read_burst_rvalid_2166 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_2166 <= 0;
            read_burst_rlast_2167 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_2166 <= 0;
            read_burst_rlast_2167 <= 0;
          end 
          if(read_burst_rlast_2167 && read_burst_rvalid_2166 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_35 <= read_burst_fsm_35_init;
          end 
          if(0) begin
            read_burst_fsm_35 <= read_burst_fsm_35_init;
          end 
        end
      endcase
    end
  end

  localparam control_matmul_16_1 = 1;
  localparam control_matmul_16_2 = 2;
  localparam control_matmul_16_3 = 3;
  localparam control_matmul_16_4 = 4;
  localparam control_matmul_16_5 = 5;
  localparam control_matmul_16_6 = 6;
  localparam control_matmul_16_7 = 7;
  localparam control_matmul_16_8 = 8;
  localparam control_matmul_16_9 = 9;
  localparam control_matmul_16_10 = 10;
  localparam control_matmul_16_11 = 11;
  localparam control_matmul_16_12 = 12;
  localparam control_matmul_16_13 = 13;
  localparam control_matmul_16_14 = 14;
  localparam control_matmul_16_15 = 15;
  localparam control_matmul_16_16 = 16;
  localparam control_matmul_16_17 = 17;
  localparam control_matmul_16_18 = 18;
  localparam control_matmul_16_19 = 19;
  localparam control_matmul_16_20 = 20;
  localparam control_matmul_16_21 = 21;
  localparam control_matmul_16_22 = 22;
  localparam control_matmul_16_23 = 23;
  localparam control_matmul_16_24 = 24;
  localparam control_matmul_16_25 = 25;
  localparam control_matmul_16_26 = 26;
  localparam control_matmul_16_27 = 27;
  localparam control_matmul_16_28 = 28;

  always @(posedge CLK) begin
    if(RST) begin
      control_matmul_16 <= control_matmul_16_init;
      _control_matmul_16_called <= 0;
      matmul_16_filter_base_offset <= 0;
      matmul_16_filter_page_comp_offset <= 0;
      matmul_16_filter_page_dma_offset <= 0;
      matmul_16_act_base_offset_row <= 0;
      matmul_16_act_base_offset_bat <= 0;
      matmul_16_dma_flag_0 <= 0;
      matmul_16_act_page_comp_offset_0 <= 0;
      matmul_16_act_page_dma_offset_0 <= 0;
      matmul_16_out_base_offset_val <= 0;
      matmul_16_out_base_offset_col <= 0;
      matmul_16_out_base_offset_row <= 0;
      matmul_16_out_base_offset_bat <= 0;
      matmul_16_out_base_offset_och <= 0;
      matmul_16_out_page <= 0;
      matmul_16_out_page_comp_offset <= 0;
      matmul_16_out_page_dma_offset <= 0;
      matmul_16_out_laddr_offset <= 0;
      matmul_16_sync_out_count <= 0;
      matmul_16_write_count <= 0;
      matmul_16_next_out_write_size <= 0;
      matmul_16_row_count <= 0;
      matmul_16_bat_count <= 0;
      matmul_16_och_count <= 0;
      matmul_16_row_select <= 0;
      matmul_16_prev_row_count <= 0;
      matmul_16_prev_bat_count <= 0;
      matmul_16_prev_och_count <= 0;
      matmul_16_prev_row_select <= 0;
      matmul_16_out_col_count <= 0;
      matmul_16_out_row_count <= 0;
      matmul_16_out_ram_select <= 0;
      matmul_16_skip_read_filter <= 0;
      matmul_16_skip_read_act <= 0;
      matmul_16_skip_comp <= 0;
      matmul_16_skip_write_out <= 1;
    end else begin
      case(control_matmul_16)
        control_matmul_16_init: begin
          if(main_fsm == 39) begin
            _control_matmul_16_called <= 1;
          end 
          if(main_fsm == 49) begin
            _control_matmul_16_called <= 1;
          end 
          if(main_fsm == 39) begin
            control_matmul_16 <= control_matmul_16_1;
          end 
          if(main_fsm == 49) begin
            control_matmul_16 <= control_matmul_16_1;
          end 
        end
        control_matmul_16_1: begin
          control_matmul_16 <= control_matmul_16_2;
        end
        control_matmul_16_2: begin
          matmul_16_filter_base_offset <= 0;
          matmul_16_filter_page_comp_offset <= 0;
          matmul_16_filter_page_dma_offset <= 0;
          matmul_16_act_base_offset_row <= 0;
          matmul_16_act_base_offset_bat <= 0;
          matmul_16_dma_flag_0 <= 1;
          matmul_16_act_page_comp_offset_0 <= 0;
          matmul_16_act_page_dma_offset_0 <= 0;
          matmul_16_out_base_offset_val <= 0;
          matmul_16_out_base_offset_col <= 0;
          matmul_16_out_base_offset_row <= 0;
          matmul_16_out_base_offset_bat <= 0;
          matmul_16_out_base_offset_och <= 0;
          matmul_16_out_page <= 0;
          matmul_16_out_page_comp_offset <= 0;
          matmul_16_out_page_dma_offset <= 0;
          matmul_16_out_laddr_offset <= 0;
          matmul_16_sync_out_count <= 0;
          matmul_16_write_count <= 0;
          matmul_16_next_out_write_size <= (cparam_matmul_16_max_och_count == 0)? cparam_matmul_16_out_write_size_res : cparam_matmul_16_out_write_size;
          matmul_16_row_count <= 0;
          matmul_16_bat_count <= 0;
          matmul_16_och_count <= 0;
          matmul_16_row_select <= 0;
          matmul_16_prev_row_count <= 0;
          matmul_16_prev_bat_count <= 0;
          matmul_16_prev_och_count <= 0;
          matmul_16_prev_row_select <= 0;
          matmul_16_out_col_count <= 0;
          matmul_16_out_row_count <= 0;
          matmul_16_out_ram_select <= 0;
          matmul_16_skip_read_filter <= 0;
          matmul_16_skip_read_act <= 0;
          matmul_16_skip_comp <= 0;
          matmul_16_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_matmul_16 <= control_matmul_16_3;
          end 
        end
        control_matmul_16_3: begin
          if(_maxi_read_idle) begin
            control_matmul_16 <= control_matmul_16_4;
          end 
        end
        control_matmul_16_4: begin
          if(_maxi_read_req_idle) begin
            control_matmul_16 <= control_matmul_16_5;
          end 
        end
        control_matmul_16_5: begin
          if(_maxi_read_idle) begin
            control_matmul_16 <= control_matmul_16_6;
          end 
        end
        control_matmul_16_6: begin
          if(cparam_matmul_16_data_stationary == 0) begin
            control_matmul_16 <= control_matmul_16_7;
          end 
          if(cparam_matmul_16_data_stationary == 1) begin
            control_matmul_16 <= control_matmul_16_12;
          end 
        end
        control_matmul_16_7: begin
          control_matmul_16 <= control_matmul_16_8;
          if(matmul_16_skip_read_filter) begin
            control_matmul_16 <= control_matmul_16_11;
          end 
        end
        control_matmul_16_8: begin
          if(_maxi_read_req_idle) begin
            control_matmul_16 <= control_matmul_16_9;
          end 
        end
        control_matmul_16_9: begin
          if(_maxi_read_idle) begin
            control_matmul_16 <= control_matmul_16_10;
          end 
        end
        control_matmul_16_10: begin
          control_matmul_16 <= control_matmul_16_11;
        end
        control_matmul_16_11: begin
          if(cparam_matmul_16_data_stationary == 0) begin
            control_matmul_16 <= control_matmul_16_12;
          end 
          if(cparam_matmul_16_data_stationary == 1) begin
            control_matmul_16 <= control_matmul_16_18;
          end 
        end
        control_matmul_16_12: begin
          control_matmul_16 <= control_matmul_16_13;
          if(matmul_16_skip_read_act) begin
            control_matmul_16 <= control_matmul_16_17;
          end 
        end
        control_matmul_16_13: begin
          control_matmul_16 <= control_matmul_16_14;
          if(matmul_16_mux_dma_pad_mask_0 || !matmul_16_mux_dma_flag_0) begin
            control_matmul_16 <= control_matmul_16_16;
          end 
        end
        control_matmul_16_14: begin
          if(_maxi_read_req_idle) begin
            control_matmul_16 <= control_matmul_16_15;
          end 
        end
        control_matmul_16_15: begin
          if(_maxi_read_idle) begin
            control_matmul_16 <= control_matmul_16_16;
          end 
        end
        control_matmul_16_16: begin
          control_matmul_16 <= control_matmul_16_17;
        end
        control_matmul_16_17: begin
          if(cparam_matmul_16_data_stationary == 0) begin
            control_matmul_16 <= control_matmul_16_18;
          end 
          if(cparam_matmul_16_data_stationary == 1) begin
            control_matmul_16 <= control_matmul_16_7;
          end 
        end
        control_matmul_16_18: begin
          if(_maxi_write_idle) begin
            control_matmul_16 <= control_matmul_16_19;
          end 
        end
        control_matmul_16_19: begin
          if(matmul_16_comp_fsm == 0) begin
            control_matmul_16 <= control_matmul_16_20;
          end 
        end
        control_matmul_16_20: begin
          control_matmul_16 <= control_matmul_16_21;
          if(matmul_16_skip_write_out) begin
            control_matmul_16 <= control_matmul_16_26;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_prev_och_count < cparam_matmul_16_max_och_count)) begin
            control_matmul_16 <= control_matmul_16_26;
          end 
        end
        control_matmul_16_21: begin
          if(matmul_16_sync_comp_count >= matmul_16_sync_out_count + cparam_matmul_16_inc_sync_out) begin
            control_matmul_16 <= control_matmul_16_22;
          end 
        end
        control_matmul_16_22: begin
          if(!matmul_16_dma_out_mask_0) begin
            control_matmul_16 <= control_matmul_16_23;
          end 
          if(matmul_16_dma_out_mask_0) begin
            control_matmul_16 <= control_matmul_16_24;
          end 
        end
        control_matmul_16_23: begin
          if(_maxi_write_req_idle) begin
            control_matmul_16 <= control_matmul_16_24;
          end 
        end
        control_matmul_16_24: begin
          control_matmul_16 <= control_matmul_16_25;
        end
        control_matmul_16_25: begin
          matmul_16_write_count <= matmul_16_write_count + 1;
          if(matmul_16_out_ram_select == 0) begin
            matmul_16_out_laddr_offset <= matmul_16_out_laddr_offset + matmul_16_next_out_write_size;
          end 
          if((cparam_matmul_16_data_stationary == 0) && !cparam_matmul_16_keep_filter) begin
            matmul_16_out_base_offset_col <= matmul_16_out_base_offset_col + cparam_matmul_16_out_col_step;
            matmul_16_out_col_count <= matmul_16_out_col_count + 1;
          end 
          matmul_16_out_ram_select <= matmul_16_out_ram_select + 1;
          if(matmul_16_out_ram_select == 0) begin
            matmul_16_out_ram_select <= 0;
          end 
          matmul_16_sync_out_count <= matmul_16_sync_out_count + cparam_matmul_16_inc_sync_out;
          if((cparam_matmul_16_data_stationary == 0) && !cparam_matmul_16_keep_filter && (matmul_16_write_count >= cparam_matmul_16_out_num_col - 1) || (cparam_matmul_16_data_stationary == 0) && cparam_matmul_16_keep_filter || (cparam_matmul_16_data_stationary == 1)) begin
            matmul_16_sync_out_count <= matmul_16_sync_out_count + (cparam_matmul_16_inc_sync_out + cparam_matmul_16_inc_sync_out_res);
          end 
          if((cparam_matmul_16_data_stationary == 0) && !cparam_matmul_16_keep_filter) begin
            control_matmul_16 <= control_matmul_16_20;
          end 
          if((cparam_matmul_16_data_stationary == 0) && !cparam_matmul_16_keep_filter && (matmul_16_write_count >= cparam_matmul_16_out_num_col - 1) || (cparam_matmul_16_data_stationary == 0) && cparam_matmul_16_keep_filter || (cparam_matmul_16_data_stationary == 1)) begin
            control_matmul_16 <= control_matmul_16_26;
          end 
        end
        control_matmul_16_26: begin
          if(matmul_16_update_filter) begin
            matmul_16_filter_base_offset <= matmul_16_filter_base_offset + cparam_matmul_16_filter_base_step;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_och_count >= cparam_matmul_16_max_och_count)) begin
            matmul_16_filter_base_offset <= 0;
          end 
          if(matmul_16_update_filter) begin
            matmul_16_och_count <= matmul_16_och_count + cparam_matmul_16_och_count_step;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_och_count >= cparam_matmul_16_max_och_count)) begin
            matmul_16_och_count <= 0;
          end 
          if(matmul_16_update_filter) begin
            matmul_16_filter_page_comp_offset <= matmul_16_filter_page_comp_offset + cparam_matmul_16_filter_read_step;
            matmul_16_filter_page_dma_offset <= matmul_16_filter_page_dma_offset + cparam_matmul_16_filter_read_step;
          end 
          if(matmul_16_update_filter && (matmul_16_filter_page_comp_offset + cparam_matmul_16_filter_read_step + cparam_matmul_16_filter_read_step > 16384)) begin
            matmul_16_filter_page_comp_offset <= 0;
            matmul_16_filter_page_dma_offset <= 0;
          end 
          if(matmul_16_update_act) begin
            matmul_16_act_base_offset_row <= matmul_16_act_base_offset_row + cparam_matmul_16_act_row_step;
          end 
          if(matmul_16_update_act && (matmul_16_row_count >= cparam_matmul_16_max_row_count)) begin
            matmul_16_act_base_offset_row <= 0;
            matmul_16_act_base_offset_bat <= matmul_16_act_base_offset_bat + cparam_matmul_16_act_bat_step;
          end 
          if(matmul_16_update_act && (matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count)) begin
            matmul_16_act_base_offset_bat <= 0;
          end 
          if(!matmul_16_update_act) begin
            matmul_16_dma_flag_0 <= 0;
          end 
          if(matmul_16_update_act) begin
            matmul_16_dma_flag_0 <= cparam_matmul_16_dma_flag_conds_0;
          end 
          if(matmul_16_update_act && (matmul_16_row_count >= cparam_matmul_16_max_row_count)) begin
            matmul_16_dma_flag_0 <= 1;
          end 
          if(matmul_16_update_act) begin
            matmul_16_row_count <= matmul_16_row_count + cparam_matmul_16_stride_row_par_row;
          end 
          if(matmul_16_update_act && (matmul_16_row_count >= cparam_matmul_16_max_row_count)) begin
            matmul_16_row_count <= 0;
            matmul_16_bat_count <= matmul_16_bat_count + 1;
          end 
          if(matmul_16_update_act && (matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count)) begin
            matmul_16_bat_count <= 0;
          end 
          if(matmul_16_update_act && (cparam_matmul_16_stride_row_par_row < 1)) begin
            matmul_16_row_select <= matmul_16_row_select + cparam_matmul_16_stride_row_par_row;
            matmul_16_prev_row_select <= matmul_16_row_select;
          end 
          if(matmul_16_update_act && (cparam_matmul_16_stride_row_par_row < 1) && (matmul_16_row_select + cparam_matmul_16_stride_row_par_row >= 1)) begin
            matmul_16_row_select <= matmul_16_row_select - (1 - cparam_matmul_16_stride_row_par_row);
            matmul_16_prev_row_select <= matmul_16_row_select;
          end 
          if(matmul_16_update_act && !(cparam_matmul_16_stride_row_par_row < 1)) begin
            matmul_16_row_select <= 0;
            matmul_16_prev_row_select <= 0;
          end 
          if(matmul_16_update_act && (matmul_16_row_count >= cparam_matmul_16_max_row_count)) begin
            matmul_16_row_select <= 0;
            matmul_16_prev_row_select <= 0;
          end 
          if(matmul_16_update_act && matmul_16_mux_next_dma_flag_0) begin
            matmul_16_act_page_comp_offset_0 <= matmul_16_act_page_comp_offset_0 + cparam_matmul_16_act_read_step;
            matmul_16_act_page_dma_offset_0 <= matmul_16_act_page_dma_offset_0 + cparam_matmul_16_act_read_step;
          end 
          if(matmul_16_update_act && matmul_16_mux_next_dma_flag_0 && (matmul_16_act_page_comp_offset_0 + cparam_matmul_16_act_read_step + cparam_matmul_16_act_read_step > 8192)) begin
            matmul_16_act_page_comp_offset_0 <= 0;
            matmul_16_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_matmul_16_data_stationary == 0) && (matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count) && cparam_matmul_16_keep_input) begin
            matmul_16_act_page_comp_offset_0 <= 0;
            matmul_16_act_page_dma_offset_0 <= 0;
          end 
          matmul_16_next_out_write_size <= (matmul_16_och_count >= cparam_matmul_16_max_och_count)? cparam_matmul_16_out_write_size_res : cparam_matmul_16_out_write_size;
          if(!matmul_16_skip_write_out) begin
            matmul_16_write_count <= 0;
            matmul_16_out_laddr_offset <= 0;
            matmul_16_out_ram_select <= 0;
          end 
          if((cparam_matmul_16_data_stationary == 0) && !matmul_16_skip_write_out) begin
            matmul_16_out_base_offset_col <= 0;
            matmul_16_out_base_offset_row <= matmul_16_out_base_offset_row + cparam_matmul_16_out_row_step;
            matmul_16_out_col_count <= 0;
            matmul_16_out_row_count <= matmul_16_out_row_count + 1;
          end 
          if((cparam_matmul_16_data_stationary == 0) && !matmul_16_skip_write_out && (matmul_16_prev_row_count >= cparam_matmul_16_max_row_count)) begin
            matmul_16_out_base_offset_row <= 0;
            matmul_16_out_base_offset_bat <= matmul_16_out_base_offset_bat + cparam_matmul_16_out_bat_step;
            matmul_16_out_row_count <= 0;
          end 
          if((cparam_matmul_16_data_stationary == 0) && !matmul_16_skip_write_out && (matmul_16_prev_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_prev_bat_count >= cparam_matmul_16_max_bat_count)) begin
            matmul_16_out_base_offset_bat <= 0;
            matmul_16_out_base_offset_och <= matmul_16_out_base_offset_och + cparam_matmul_16_out_och_step;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_prev_och_count >= cparam_matmul_16_max_och_count) && !matmul_16_skip_write_out) begin
            matmul_16_out_base_offset_row <= matmul_16_out_base_offset_row + cparam_matmul_16_out_row_step;
          end 
          if((cparam_matmul_16_data_stationary == 0) && !matmul_16_out_page) begin
            matmul_16_out_page_comp_offset <= 64;
            matmul_16_out_page_dma_offset <= 0;
            matmul_16_out_page <= 1;
          end 
          if((cparam_matmul_16_data_stationary == 0) && matmul_16_out_page) begin
            matmul_16_out_page_comp_offset <= 0;
            matmul_16_out_page_dma_offset <= 64;
            matmul_16_out_page <= 0;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_och_count >= cparam_matmul_16_max_och_count) && !matmul_16_out_page) begin
            matmul_16_out_page_comp_offset <= 64;
            matmul_16_out_page_dma_offset <= 0;
            matmul_16_out_page <= 1;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_och_count >= cparam_matmul_16_max_och_count) && matmul_16_out_page) begin
            matmul_16_out_page_comp_offset <= 0;
            matmul_16_out_page_dma_offset <= 64;
            matmul_16_out_page <= 0;
          end 
          matmul_16_prev_row_count <= matmul_16_row_count;
          matmul_16_prev_bat_count <= matmul_16_bat_count;
          matmul_16_prev_och_count <= matmul_16_och_count;
          if((matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count) && (matmul_16_och_count >= cparam_matmul_16_max_och_count)) begin
            matmul_16_skip_read_filter <= 1;
          end 
          if((cparam_matmul_16_data_stationary == 1) && cparam_matmul_16_keep_filter) begin
            matmul_16_skip_read_filter <= 1;
          end 
          if((matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count) && (matmul_16_och_count >= cparam_matmul_16_max_och_count)) begin
            matmul_16_skip_read_act <= 1;
          end 
          if((cparam_matmul_16_data_stationary == 0) && (matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count) && cparam_matmul_16_keep_input) begin
            matmul_16_skip_read_act <= 1;
          end 
          if((matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count) && (matmul_16_och_count >= cparam_matmul_16_max_och_count)) begin
            matmul_16_skip_comp <= 1;
          end 
          if(matmul_16_skip_write_out && (matmul_16_prev_row_count == 0) && (matmul_16_prev_bat_count == 0) && (matmul_16_prev_och_count == 0)) begin
            matmul_16_skip_write_out <= 0;
          end 
          if(cparam_matmul_16_data_stationary == 0) begin
            control_matmul_16 <= control_matmul_16_12;
          end 
          if((cparam_matmul_16_data_stationary == 0) && (matmul_16_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_bat_count >= cparam_matmul_16_max_bat_count)) begin
            control_matmul_16 <= control_matmul_16_7;
          end 
          if(cparam_matmul_16_data_stationary == 1) begin
            control_matmul_16 <= control_matmul_16_7;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_och_count >= cparam_matmul_16_max_och_count)) begin
            control_matmul_16 <= control_matmul_16_12;
          end 
          if(!matmul_16_skip_write_out && (matmul_16_prev_och_count >= cparam_matmul_16_max_och_count) && (matmul_16_prev_row_count >= cparam_matmul_16_max_row_count) && (matmul_16_prev_bat_count >= cparam_matmul_16_max_bat_count)) begin
            control_matmul_16 <= control_matmul_16_27;
          end 
        end
        control_matmul_16_27: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_matmul_16 <= control_matmul_16_28;
          end 
        end
        control_matmul_16_28: begin
          if(main_fsm == 42) begin
            _control_matmul_16_called <= 0;
          end 
          if(main_fsm == 52) begin
            _control_matmul_16_called <= 0;
          end 
          if(main_fsm == 42) begin
            control_matmul_16 <= control_matmul_16_init;
          end 
          if(main_fsm == 52) begin
            control_matmul_16 <= control_matmul_16_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_36_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_36 <= write_burst_fsm_36_init;
      write_burst_addr_2173 <= 0;
      write_burst_stride_2174 <= 0;
      write_burst_length_2175 <= 0;
      write_burst_done_2176 <= 0;
    end else begin
      case(write_burst_fsm_36)
        write_burst_fsm_36_init: begin
          write_burst_addr_2173 <= _maxi_read_local_addr_buf;
          write_burst_stride_2174 <= _maxi_read_local_stride_buf;
          write_burst_length_2175 <= _maxi_read_local_size_buf;
          write_burst_done_2176 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 8) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_36 <= write_burst_fsm_36_1;
          end 
        end
        write_burst_fsm_36_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_2173 <= write_burst_addr_2173 + write_burst_stride_2174;
            write_burst_length_2175 <= write_burst_length_2175 - 1;
            write_burst_done_2176 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2175 <= 1)) begin
            write_burst_done_2176 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_2176 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2175 <= 1)) begin
            write_burst_fsm_36 <= write_burst_fsm_36_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_36 <= write_burst_fsm_36_init;
          end 
          if(0) begin
            write_burst_fsm_36 <= write_burst_fsm_36_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_37_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_37 <= write_burst_fsm_37_init;
      write_burst_addr_2179 <= 0;
      write_burst_stride_2180 <= 0;
      write_burst_length_2181 <= 0;
      write_burst_done_2182 <= 0;
    end else begin
      case(write_burst_fsm_37)
        write_burst_fsm_37_init: begin
          write_burst_addr_2179 <= _maxi_read_local_addr_buf;
          write_burst_stride_2180 <= _maxi_read_local_stride_buf;
          write_burst_length_2181 <= _maxi_read_local_size_buf;
          write_burst_done_2182 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 9) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_37 <= write_burst_fsm_37_1;
          end 
        end
        write_burst_fsm_37_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_2179 <= write_burst_addr_2179 + write_burst_stride_2180;
            write_burst_length_2181 <= write_burst_length_2181 - 1;
            write_burst_done_2182 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2181 <= 1)) begin
            write_burst_done_2182 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_2182 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2181 <= 1)) begin
            write_burst_fsm_37 <= write_burst_fsm_37_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_37 <= write_burst_fsm_37_init;
          end 
          if(0) begin
            write_burst_fsm_37 <= write_burst_fsm_37_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_38_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_38 <= write_burst_fsm_38_init;
      write_burst_addr_2187 <= 0;
      write_burst_stride_2188 <= 0;
      write_burst_length_2189 <= 0;
      write_burst_done_2190 <= 0;
    end else begin
      case(write_burst_fsm_38)
        write_burst_fsm_38_init: begin
          write_burst_addr_2187 <= _maxi_read_local_addr_buf;
          write_burst_stride_2188 <= _maxi_read_local_stride_buf;
          write_burst_length_2189 <= _maxi_read_local_size_buf;
          write_burst_done_2190 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 10) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_38 <= write_burst_fsm_38_1;
          end 
        end
        write_burst_fsm_38_1: begin
          if(write_burst_block_ram_wvalid_2185) begin
            write_burst_addr_2187 <= write_burst_addr_2187 + write_burst_stride_2188;
            write_burst_length_2189 <= write_burst_length_2189 - 1;
            write_burst_done_2190 <= 0;
          end 
          if(write_burst_block_ram_wvalid_2185 && (write_burst_length_2189 <= 1)) begin
            write_burst_done_2190 <= 1;
          end 
          if(write_burst_block_ram_wvalid_2185 && 0) begin
            write_burst_done_2190 <= 1;
          end 
          if(write_burst_block_ram_wvalid_2185 && (write_burst_length_2189 <= 1)) begin
            write_burst_fsm_38 <= write_burst_fsm_38_init;
          end 
          if(write_burst_block_ram_wvalid_2185 && 0) begin
            write_burst_fsm_38 <= write_burst_fsm_38_init;
          end 
          if(write_burst_block_ram_wquit_2186) begin
            write_burst_fsm_38 <= write_burst_fsm_38_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_39_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_39 <= write_burst_fsm_39_init;
      write_burst_addr_2193 <= 0;
      write_burst_stride_2194 <= 0;
      write_burst_length_2195 <= 0;
      write_burst_done_2196 <= 0;
    end else begin
      case(write_burst_fsm_39)
        write_burst_fsm_39_init: begin
          write_burst_addr_2193 <= _maxi_read_local_addr_buf;
          write_burst_stride_2194 <= _maxi_read_local_stride_buf;
          write_burst_length_2195 <= _maxi_read_local_size_buf;
          write_burst_done_2196 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 10) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_39 <= write_burst_fsm_39_1;
          end 
        end
        write_burst_fsm_39_1: begin
          if(write_burst_block_ram_wvalid_2191) begin
            write_burst_addr_2193 <= write_burst_addr_2193 + write_burst_stride_2194;
            write_burst_length_2195 <= write_burst_length_2195 - 1;
            write_burst_done_2196 <= 0;
          end 
          if(write_burst_block_ram_wvalid_2191 && (write_burst_length_2195 <= 1)) begin
            write_burst_done_2196 <= 1;
          end 
          if(write_burst_block_ram_wvalid_2191 && 0) begin
            write_burst_done_2196 <= 1;
          end 
          if(write_burst_block_ram_wvalid_2191 && (write_burst_length_2195 <= 1)) begin
            write_burst_fsm_39 <= write_burst_fsm_39_init;
          end 
          if(write_burst_block_ram_wvalid_2191 && 0) begin
            write_burst_fsm_39 <= write_burst_fsm_39_init;
          end 
          if(write_burst_block_ram_wquit_2192) begin
            write_burst_fsm_39 <= write_burst_fsm_39_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_40_1 = 1;
  localparam write_burst_block_fsm_40_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_40 <= write_burst_block_fsm_40_init;
      write_burst_block_length_2197 <= 0;
      write_burst_block_blocksize_2198 <= 0;
      write_burst_block_done_2199 <= 0;
      write_burst_block_count_2200 <= 0;
    end else begin
      case(write_burst_block_fsm_40)
        write_burst_block_fsm_40_init: begin
          write_burst_block_length_2197 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_2198 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_2199 <= 0;
          write_burst_block_count_2200 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 10) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_1;
          end 
        end
        write_burst_block_fsm_40_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_2197 <= write_burst_block_length_2197 - 1;
            write_burst_block_done_2199 <= 0;
            write_burst_block_count_2200 <= write_burst_block_count_2200 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_2197 <= 1)) begin
            write_burst_block_done_2199 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_2199 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_2200 == write_burst_block_blocksize_2198 - 1)) begin
            write_burst_block_count_2200 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_2200 == write_burst_block_blocksize_2198 - 1)) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_2197 <= 1)) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_init;
          end 
          if(0) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_init;
          end 
        end
        write_burst_block_fsm_40_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_2197 <= write_burst_block_length_2197 - 1;
            write_burst_block_done_2199 <= 0;
            write_burst_block_count_2200 <= write_burst_block_count_2200 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_2197 <= 1)) begin
            write_burst_block_done_2199 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_2199 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_2200 == write_burst_block_blocksize_2198 - 1)) begin
            write_burst_block_count_2200 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_2200 == write_burst_block_blocksize_2198 - 1)) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_2197 <= 1)) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_init;
          end 
          if(0) begin
            write_burst_block_fsm_40 <= write_burst_block_fsm_40_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_41_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_41 <= write_burst_fsm_41_init;
      write_burst_addr_2203 <= 0;
      write_burst_stride_2204 <= 0;
      write_burst_length_2205 <= 0;
      write_burst_done_2206 <= 0;
    end else begin
      case(write_burst_fsm_41)
        write_burst_fsm_41_init: begin
          write_burst_addr_2203 <= _maxi_read_local_addr_buf;
          write_burst_stride_2204 <= _maxi_read_local_stride_buf;
          write_burst_length_2205 <= _maxi_read_local_size_buf;
          write_burst_done_2206 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 11) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_41 <= write_burst_fsm_41_1;
          end 
        end
        write_burst_fsm_41_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_2203 <= write_burst_addr_2203 + write_burst_stride_2204;
            write_burst_length_2205 <= write_burst_length_2205 - 1;
            write_burst_done_2206 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2205 <= 1)) begin
            write_burst_done_2206 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_2206 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_2205 <= 1)) begin
            write_burst_fsm_41 <= write_burst_fsm_41_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_41 <= write_burst_fsm_41_init;
          end 
          if(0) begin
            write_burst_fsm_41 <= write_burst_fsm_41_init;
          end 
        end
      endcase
    end
  end

  localparam matmul_16_comp_fsm_1 = 1;
  localparam matmul_16_comp_fsm_2 = 2;
  localparam matmul_16_comp_fsm_3 = 3;
  localparam matmul_16_comp_fsm_4 = 4;
  localparam matmul_16_comp_fsm_5 = 5;
  localparam matmul_16_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      matmul_16_comp_fsm <= matmul_16_comp_fsm_init;
      matmul_16_stream_act_local_0 <= 0;
      matmul_16_stream_out_local_col <= 0;
      matmul_16_stream_out_local_val <= 0;
      matmul_16_col_count <= 0;
      matmul_16_col_select <= 0;
      matmul_16_filter_page_comp_offset_buf <= 0;
      matmul_16_act_page_comp_offset_buf_0 <= 0;
      matmul_16_out_page_comp_offset_buf <= 0;
      matmul_16_row_count_buf <= 0;
      matmul_16_row_select_buf <= 0;
      matmul_16_och_count_buf <= 0;
      matmul_16_next_stream_num_ops <= 0;
      matmul_16_stream_pad_masks <= 0;
      matmul_16_sync_comp_count <= 0;
    end else begin
      if(_stream_matmul_16_sink_stop) begin
        matmul_16_sync_comp_count <= matmul_16_sync_comp_count + 1;
      end 
      if(control_matmul_16 == 6) begin
        matmul_16_sync_comp_count <= 0;
      end 
      case(matmul_16_comp_fsm)
        matmul_16_comp_fsm_init: begin
          if((control_matmul_16 == 19) && !matmul_16_skip_comp) begin
            matmul_16_comp_fsm <= matmul_16_comp_fsm_1;
          end 
        end
        matmul_16_comp_fsm_1: begin
          matmul_16_stream_act_local_0 <= 0;
          if(cparam_matmul_16_stream_act_local_small_flags_0) begin
            matmul_16_stream_act_local_0 <= cparam_matmul_16_stream_act_local_small_offset;
          end 
          if(cparam_matmul_16_stream_act_local_large_flags_0) begin
            matmul_16_stream_act_local_0 <= cparam_matmul_16_stream_act_local_large_offset;
          end 
          matmul_16_stream_out_local_col <= 0;
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_och_count == 0)) begin
            matmul_16_stream_out_local_val <= 0;
          end 
          matmul_16_col_count <= 0;
          matmul_16_col_select <= cparam_matmul_16_col_select_initval;
          matmul_16_filter_page_comp_offset_buf <= matmul_16_filter_page_comp_offset;
          matmul_16_act_page_comp_offset_buf_0 <= matmul_16_act_page_comp_offset_0;
          matmul_16_out_page_comp_offset_buf <= matmul_16_out_page_comp_offset;
          matmul_16_row_count_buf <= matmul_16_row_count;
          matmul_16_row_select_buf <= matmul_16_row_select;
          matmul_16_och_count_buf <= matmul_16_och_count;
          matmul_16_next_stream_num_ops <= (matmul_16_och_count >= cparam_matmul_16_max_och_count)? cparam_matmul_16_stream_num_ops_res : cparam_matmul_16_stream_num_ops;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_2;
        end
        matmul_16_comp_fsm_2: begin
          matmul_16_stream_pad_masks <= { matmul_16_stream_pad_mask_0_0 };
          matmul_16_comp_fsm <= matmul_16_comp_fsm_3;
        end
        matmul_16_comp_fsm_3: begin
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          if(_stream_matmul_16_stream_oready) begin
            matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
          end 
          matmul_16_comp_fsm <= matmul_16_comp_fsm_4;
        end
        matmul_16_comp_fsm_4: begin
          if(!_stream_matmul_16_source_busy) begin
            matmul_16_comp_fsm <= matmul_16_comp_fsm_5;
          end 
        end
        matmul_16_comp_fsm_5: begin
          if(_stream_matmul_16_busy) begin
            matmul_16_comp_fsm <= matmul_16_comp_fsm_6;
          end 
        end
        matmul_16_comp_fsm_6: begin
          if(!((matmul_16_col_select == 0)? cparam_matmul_16_inc_act_laddr_conds_0 : 0)) begin
            matmul_16_stream_act_local_0 <= matmul_16_stream_act_local_0 + cparam_matmul_16_inc_act_laddr_small;
          end 
          if((matmul_16_col_select == 0)? cparam_matmul_16_inc_act_laddr_conds_0 : 0) begin
            matmul_16_stream_act_local_0 <= matmul_16_stream_act_local_0 + cparam_matmul_16_inc_act_laddr_large;
          end 
          if(matmul_16_col_count >= cparam_matmul_16_max_col_count) begin
            matmul_16_stream_act_local_0 <= 0;
          end 
          if((matmul_16_col_count >= cparam_matmul_16_max_col_count) && cparam_matmul_16_stream_act_local_small_flags_0) begin
            matmul_16_stream_act_local_0 <= cparam_matmul_16_stream_act_local_small_offset;
          end 
          if((matmul_16_col_count >= cparam_matmul_16_max_col_count) && cparam_matmul_16_stream_act_local_large_flags_0) begin
            matmul_16_stream_act_local_0 <= cparam_matmul_16_stream_act_local_large_offset;
          end 
          if(cparam_matmul_16_data_stationary == 0) begin
            matmul_16_stream_out_local_col <= matmul_16_stream_out_local_col + matmul_16_next_stream_num_ops;
          end 
          if((cparam_matmul_16_data_stationary == 0) && (matmul_16_col_count >= cparam_matmul_16_max_col_count)) begin
            matmul_16_stream_out_local_col <= 0;
          end 
          if(cparam_matmul_16_data_stationary == 1) begin
            matmul_16_stream_out_local_col <= matmul_16_stream_out_local_col + cparam_matmul_16_inc_out_laddr_col;
          end 
          if((cparam_matmul_16_data_stationary == 1) && (matmul_16_col_count >= cparam_matmul_16_max_col_count)) begin
            matmul_16_stream_out_local_val <= matmul_16_stream_out_local_val + matmul_16_next_stream_num_ops;
            matmul_16_stream_out_local_col <= 0;
          end 
          matmul_16_col_count <= matmul_16_col_count + cparam_matmul_16_stride_col_par_col;
          if(matmul_16_col_count >= cparam_matmul_16_max_col_count) begin
            matmul_16_col_count <= 0;
          end 
          matmul_16_col_select <= matmul_16_col_select + cparam_matmul_16_stride_col_mod_filter_num;
          if(matmul_16_col_select + cparam_matmul_16_stride_col_mod_filter_num >= 1) begin
            matmul_16_col_select <= matmul_16_col_select - cparam_matmul_16_filter_num_col_minus_stride_col_mod;
          end 
          if(matmul_16_col_count >= cparam_matmul_16_max_col_count) begin
            matmul_16_col_select <= cparam_matmul_16_col_select_initval;
          end 
          matmul_16_comp_fsm <= matmul_16_comp_fsm_2;
          if(matmul_16_col_count >= cparam_matmul_16_max_col_count) begin
            matmul_16_comp_fsm <= matmul_16_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_16_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_matmul_16_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_source_7_source_pat_fsm_0 <= _stream_matmul_16_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_matmul_16_source_7_source_pat_fsm_0)
        _stream_matmul_16_source_7_source_pat_fsm_0_init: begin
          if(_stream_matmul_16_source_start && _stream_matmul_16_source_7_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_7_source_pat_fsm_0 <= _stream_matmul_16_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_matmul_16_source_7_source_pat_fsm_0_1: begin
          if(_stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_7_source_pat_fsm_0 <= _stream_matmul_16_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_matmul_16_source_7_pat_count_0 == 0) && (_source_stream_matmul_16_source_7_pat_count_1 == 0) && (_source_stream_matmul_16_source_7_pat_count_2 == 0) && (_source_stream_matmul_16_source_7_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_7_source_pat_fsm_0 <= _stream_matmul_16_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_matmul_16_source_7_source_pat_fsm_0_2: begin
          if(_stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_7_source_pat_fsm_0 <= _stream_matmul_16_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_16_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_matmul_16_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_source_9_source_pat_fsm_1 <= _stream_matmul_16_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_matmul_16_source_9_source_pat_fsm_1)
        _stream_matmul_16_source_9_source_pat_fsm_1_init: begin
          if(_stream_matmul_16_source_start && _stream_matmul_16_source_9_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_9_source_pat_fsm_1 <= _stream_matmul_16_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_matmul_16_source_9_source_pat_fsm_1_1: begin
          if(_stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_9_source_pat_fsm_1 <= _stream_matmul_16_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_matmul_16_source_9_pat_count_0 == 0) && (_source_stream_matmul_16_source_9_pat_count_1 == 0) && (_source_stream_matmul_16_source_9_pat_count_2 == 0) && (_source_stream_matmul_16_source_9_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_9_source_pat_fsm_1 <= _stream_matmul_16_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_matmul_16_source_9_source_pat_fsm_1_2: begin
          if(_stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_9_source_pat_fsm_1 <= _stream_matmul_16_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_16_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_matmul_16_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_source_20_source_pat_fsm_2 <= _stream_matmul_16_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_matmul_16_source_20_source_pat_fsm_2)
        _stream_matmul_16_source_20_source_pat_fsm_2_init: begin
          if(_stream_matmul_16_source_start && _stream_matmul_16_source_20_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_20_source_pat_fsm_2 <= _stream_matmul_16_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_matmul_16_source_20_source_pat_fsm_2_1: begin
          if(_stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_20_source_pat_fsm_2 <= _stream_matmul_16_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_matmul_16_source_20_pat_count_0 == 0) && (_source_stream_matmul_16_source_20_pat_count_1 == 0) && (_source_stream_matmul_16_source_20_pat_count_2 == 0) && (_source_stream_matmul_16_source_20_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_20_source_pat_fsm_2 <= _stream_matmul_16_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_matmul_16_source_20_source_pat_fsm_2_2: begin
          if(_stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_20_source_pat_fsm_2 <= _stream_matmul_16_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_16_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_matmul_16_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_source_21_source_pat_fsm_3 <= _stream_matmul_16_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_matmul_16_source_21_source_pat_fsm_3)
        _stream_matmul_16_source_21_source_pat_fsm_3_init: begin
          if(_stream_matmul_16_source_start && _stream_matmul_16_source_21_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_21_source_pat_fsm_3 <= _stream_matmul_16_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_matmul_16_source_21_source_pat_fsm_3_1: begin
          if(_stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_21_source_pat_fsm_3 <= _stream_matmul_16_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_matmul_16_source_21_pat_count_0 == 0) && (_source_stream_matmul_16_source_21_pat_count_1 == 0) && (_source_stream_matmul_16_source_21_pat_count_2 == 0) && (_source_stream_matmul_16_source_21_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_21_source_pat_fsm_3 <= _stream_matmul_16_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_matmul_16_source_21_source_pat_fsm_3_2: begin
          if(_stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_21_source_pat_fsm_3 <= _stream_matmul_16_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_16_source_22_source_pat_fsm_4_1 = 1;
  localparam _stream_matmul_16_source_22_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_source_22_source_pat_fsm_4 <= _stream_matmul_16_source_22_source_pat_fsm_4_init;
    end else begin
      case(_stream_matmul_16_source_22_source_pat_fsm_4)
        _stream_matmul_16_source_22_source_pat_fsm_4_init: begin
          if(_stream_matmul_16_source_start && _stream_matmul_16_source_22_source_mode & 5'b10 && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_22_source_pat_fsm_4 <= _stream_matmul_16_source_22_source_pat_fsm_4_1;
          end 
        end
        _stream_matmul_16_source_22_source_pat_fsm_4_1: begin
          if(_stream_matmul_16_source_stop && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_22_source_pat_fsm_4 <= _stream_matmul_16_source_22_source_pat_fsm_4_init;
          end 
          if((_source_stream_matmul_16_source_22_pat_count_0 == 0) && (_source_stream_matmul_16_source_22_pat_count_1 == 0) && (_source_stream_matmul_16_source_22_pat_count_2 == 0) && (_source_stream_matmul_16_source_22_pat_count_3 == 0) && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_22_source_pat_fsm_4 <= _stream_matmul_16_source_22_source_pat_fsm_4_2;
          end 
        end
        _stream_matmul_16_source_22_source_pat_fsm_4_2: begin
          if(_stream_matmul_16_stream_oready) begin
            _stream_matmul_16_source_22_source_pat_fsm_4 <= _stream_matmul_16_source_22_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_16_sink_33_sink_fsm_5_1 = 1;
  localparam _stream_matmul_16_sink_33_sink_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_16_sink_33_sink_fsm_5 <= _stream_matmul_16_sink_33_sink_fsm_5_init;
    end else begin
      case(_stream_matmul_16_sink_33_sink_fsm_5)
        _stream_matmul_16_sink_33_sink_fsm_5_init: begin
          if(_stream_matmul_16_sink_start && _stream_matmul_16_sink_33_sink_mode & 5'b1 && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_sink_33_sink_fsm_5 <= _stream_matmul_16_sink_33_sink_fsm_5_1;
          end 
        end
        _stream_matmul_16_sink_33_sink_fsm_5_1: begin
          if(_stream_matmul_16_stream_oready) begin
            _stream_matmul_16_sink_33_sink_fsm_5 <= _stream_matmul_16_sink_33_sink_fsm_5_2;
          end 
        end
        _stream_matmul_16_sink_33_sink_fsm_5_2: begin
          if(stream_matmul_16_sink_34_data && (_stream_matmul_16_sink_33_sink_count == 1) && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_sink_33_sink_fsm_5 <= _stream_matmul_16_sink_33_sink_fsm_5_init;
          end 
          if(_stream_matmul_16_sink_stop && _stream_matmul_16_stream_oready) begin
            _stream_matmul_16_sink_33_sink_fsm_5 <= _stream_matmul_16_sink_33_sink_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_42_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_42 <= read_burst_fsm_42_init;
      read_burst_addr_2492 <= 0;
      read_burst_stride_2493 <= 0;
      read_burst_length_2494 <= 0;
      read_burst_rvalid_2495 <= 0;
      read_burst_rlast_2496 <= 0;
    end else begin
      case(read_burst_fsm_42)
        read_burst_fsm_42_init: begin
          read_burst_addr_2492 <= _maxi_write_local_addr_buf;
          read_burst_stride_2493 <= _maxi_write_local_stride_buf;
          read_burst_length_2494 <= _maxi_write_size_buf;
          read_burst_rvalid_2495 <= 0;
          read_burst_rlast_2496 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 3) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_42 <= read_burst_fsm_42_1;
          end 
        end
        read_burst_fsm_42_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2494 > 0)) begin
            read_burst_addr_2492 <= read_burst_addr_2492 + read_burst_stride_2493;
            read_burst_length_2494 <= read_burst_length_2494 - 1;
            read_burst_rvalid_2495 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_2494 <= 1)) begin
            read_burst_rlast_2496 <= 1;
          end 
          if(read_burst_rlast_2496 && read_burst_rvalid_2495 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_2495 <= 0;
            read_burst_rlast_2496 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_2495 <= 0;
            read_burst_rlast_2496 <= 0;
          end 
          if(read_burst_rlast_2496 && read_burst_rvalid_2495 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_42 <= read_burst_fsm_42_init;
          end 
          if(0) begin
            read_burst_fsm_42 <= read_burst_fsm_42_init;
          end 
        end
      endcase
    end
  end


endmodule



module _maxi_read_req_fifo
(
  input CLK,
  input RST,
  input _maxi_read_req_fifo_enq,
  input [137-1:0] _maxi_read_req_fifo_wdata,
  output _maxi_read_req_fifo_full,
  output _maxi_read_req_fifo_almost_full,
  input _maxi_read_req_fifo_deq,
  output [137-1:0] _maxi_read_req_fifo_rdata,
  output _maxi_read_req_fifo_empty,
  output _maxi_read_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_read_req_fifo_full = is_full;
  assign _maxi_read_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_read_req_fifo_empty = is_empty;
  assign _maxi_read_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_read_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_read_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_read_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _maxi_write_req_fifo
(
  input CLK,
  input RST,
  input _maxi_write_req_fifo_enq,
  input [137-1:0] _maxi_write_req_fifo_wdata,
  output _maxi_write_req_fifo_full,
  output _maxi_write_req_fifo_almost_full,
  input _maxi_write_req_fifo_deq,
  output [137-1:0] _maxi_write_req_fifo_rdata,
  output _maxi_write_req_fifo_empty,
  output _maxi_write_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_write_req_fifo_full = is_full;
  assign _maxi_write_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_write_req_fifo_empty = is_empty;
  assign _maxi_write_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_write_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_write_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_write_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module ram_w32_l16384_id0
(
  input CLK,
  input [14-1:0] ram_w32_l16384_id0_0_addr,
  output [32-1:0] ram_w32_l16384_id0_0_rdata,
  input [32-1:0] ram_w32_l16384_id0_0_wdata,
  input ram_w32_l16384_id0_0_wenable,
  input ram_w32_l16384_id0_0_enable,
  input [14-1:0] ram_w32_l16384_id0_1_addr,
  output [32-1:0] ram_w32_l16384_id0_1_rdata,
  input [32-1:0] ram_w32_l16384_id0_1_wdata,
  input ram_w32_l16384_id0_1_wenable,
  input ram_w32_l16384_id0_1_enable
);

  reg [32-1:0] ram_w32_l16384_id0_0_rdata_out;
  assign ram_w32_l16384_id0_0_rdata = ram_w32_l16384_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l16384_id0_1_rdata_out;
  assign ram_w32_l16384_id0_1_rdata = ram_w32_l16384_id0_1_rdata_out;
  reg [32-1:0] mem [0:16384-1];

  always @(posedge CLK) begin
    if(ram_w32_l16384_id0_0_enable) begin
      if(ram_w32_l16384_id0_0_wenable) begin
        mem[ram_w32_l16384_id0_0_addr] <= ram_w32_l16384_id0_0_wdata;
        ram_w32_l16384_id0_0_rdata_out <= ram_w32_l16384_id0_0_wdata;
      end else begin
        ram_w32_l16384_id0_0_rdata_out <= mem[ram_w32_l16384_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l16384_id0_1_enable) begin
      if(ram_w32_l16384_id0_1_wenable) begin
        mem[ram_w32_l16384_id0_1_addr] <= ram_w32_l16384_id0_1_wdata;
        ram_w32_l16384_id0_1_rdata_out <= ram_w32_l16384_id0_1_wdata;
      end else begin
        ram_w32_l16384_id0_1_rdata_out <= mem[ram_w32_l16384_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l16384_id1
(
  input CLK,
  input [14-1:0] ram_w32_l16384_id1_0_addr,
  output [32-1:0] ram_w32_l16384_id1_0_rdata,
  input [32-1:0] ram_w32_l16384_id1_0_wdata,
  input ram_w32_l16384_id1_0_wenable,
  input ram_w32_l16384_id1_0_enable,
  input [14-1:0] ram_w32_l16384_id1_1_addr,
  output [32-1:0] ram_w32_l16384_id1_1_rdata,
  input [32-1:0] ram_w32_l16384_id1_1_wdata,
  input ram_w32_l16384_id1_1_wenable,
  input ram_w32_l16384_id1_1_enable
);

  reg [32-1:0] ram_w32_l16384_id1_0_rdata_out;
  assign ram_w32_l16384_id1_0_rdata = ram_w32_l16384_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l16384_id1_1_rdata_out;
  assign ram_w32_l16384_id1_1_rdata = ram_w32_l16384_id1_1_rdata_out;
  reg [32-1:0] mem [0:16384-1];

  always @(posedge CLK) begin
    if(ram_w32_l16384_id1_0_enable) begin
      if(ram_w32_l16384_id1_0_wenable) begin
        mem[ram_w32_l16384_id1_0_addr] <= ram_w32_l16384_id1_0_wdata;
        ram_w32_l16384_id1_0_rdata_out <= ram_w32_l16384_id1_0_wdata;
      end else begin
        ram_w32_l16384_id1_0_rdata_out <= mem[ram_w32_l16384_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l16384_id1_1_enable) begin
      if(ram_w32_l16384_id1_1_wenable) begin
        mem[ram_w32_l16384_id1_1_addr] <= ram_w32_l16384_id1_1_wdata;
        ram_w32_l16384_id1_1_rdata_out <= ram_w32_l16384_id1_1_wdata;
      end else begin
        ram_w32_l16384_id1_1_rdata_out <= mem[ram_w32_l16384_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l8192_id0
(
  input CLK,
  input [13-1:0] ram_w32_l8192_id0_0_addr,
  output [32-1:0] ram_w32_l8192_id0_0_rdata,
  input [32-1:0] ram_w32_l8192_id0_0_wdata,
  input ram_w32_l8192_id0_0_wenable,
  input ram_w32_l8192_id0_0_enable,
  input [13-1:0] ram_w32_l8192_id0_1_addr,
  output [32-1:0] ram_w32_l8192_id0_1_rdata,
  input [32-1:0] ram_w32_l8192_id0_1_wdata,
  input ram_w32_l8192_id0_1_wenable,
  input ram_w32_l8192_id0_1_enable
);

  reg [32-1:0] ram_w32_l8192_id0_0_rdata_out;
  assign ram_w32_l8192_id0_0_rdata = ram_w32_l8192_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l8192_id0_1_rdata_out;
  assign ram_w32_l8192_id0_1_rdata = ram_w32_l8192_id0_1_rdata_out;
  reg [32-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w32_l8192_id0_0_enable) begin
      if(ram_w32_l8192_id0_0_wenable) begin
        mem[ram_w32_l8192_id0_0_addr] <= ram_w32_l8192_id0_0_wdata;
        ram_w32_l8192_id0_0_rdata_out <= ram_w32_l8192_id0_0_wdata;
      end else begin
        ram_w32_l8192_id0_0_rdata_out <= mem[ram_w32_l8192_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l8192_id0_1_enable) begin
      if(ram_w32_l8192_id0_1_wenable) begin
        mem[ram_w32_l8192_id0_1_addr] <= ram_w32_l8192_id0_1_wdata;
        ram_w32_l8192_id0_1_rdata_out <= ram_w32_l8192_id0_1_wdata;
      end else begin
        ram_w32_l8192_id0_1_rdata_out <= mem[ram_w32_l8192_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id0
(
  input CLK,
  input [9-1:0] ram_w32_l512_id0_0_addr,
  output [32-1:0] ram_w32_l512_id0_0_rdata,
  input [32-1:0] ram_w32_l512_id0_0_wdata,
  input ram_w32_l512_id0_0_wenable,
  input ram_w32_l512_id0_0_enable,
  input [9-1:0] ram_w32_l512_id0_1_addr,
  output [32-1:0] ram_w32_l512_id0_1_rdata,
  input [32-1:0] ram_w32_l512_id0_1_wdata,
  input ram_w32_l512_id0_1_wenable,
  input ram_w32_l512_id0_1_enable
);

  reg [32-1:0] ram_w32_l512_id0_0_rdata_out;
  assign ram_w32_l512_id0_0_rdata = ram_w32_l512_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id0_1_rdata_out;
  assign ram_w32_l512_id0_1_rdata = ram_w32_l512_id0_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id0_0_enable) begin
      if(ram_w32_l512_id0_0_wenable) begin
        mem[ram_w32_l512_id0_0_addr] <= ram_w32_l512_id0_0_wdata;
        ram_w32_l512_id0_0_rdata_out <= ram_w32_l512_id0_0_wdata;
      end else begin
        ram_w32_l512_id0_0_rdata_out <= mem[ram_w32_l512_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id0_1_enable) begin
      if(ram_w32_l512_id0_1_wenable) begin
        mem[ram_w32_l512_id0_1_addr] <= ram_w32_l512_id0_1_wdata;
        ram_w32_l512_id0_1_rdata_out <= ram_w32_l512_id0_1_wdata;
      end else begin
        ram_w32_l512_id0_1_rdata_out <= mem[ram_w32_l512_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id1
(
  input CLK,
  input [9-1:0] ram_w32_l512_id1_0_addr,
  output [32-1:0] ram_w32_l512_id1_0_rdata,
  input [32-1:0] ram_w32_l512_id1_0_wdata,
  input ram_w32_l512_id1_0_wenable,
  input ram_w32_l512_id1_0_enable,
  input [9-1:0] ram_w32_l512_id1_1_addr,
  output [32-1:0] ram_w32_l512_id1_1_rdata,
  input [32-1:0] ram_w32_l512_id1_1_wdata,
  input ram_w32_l512_id1_1_wenable,
  input ram_w32_l512_id1_1_enable
);

  reg [32-1:0] ram_w32_l512_id1_0_rdata_out;
  assign ram_w32_l512_id1_0_rdata = ram_w32_l512_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id1_1_rdata_out;
  assign ram_w32_l512_id1_1_rdata = ram_w32_l512_id1_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id1_0_enable) begin
      if(ram_w32_l512_id1_0_wenable) begin
        mem[ram_w32_l512_id1_0_addr] <= ram_w32_l512_id1_0_wdata;
        ram_w32_l512_id1_0_rdata_out <= ram_w32_l512_id1_0_wdata;
      end else begin
        ram_w32_l512_id1_0_rdata_out <= mem[ram_w32_l512_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id1_1_enable) begin
      if(ram_w32_l512_id1_1_wenable) begin
        mem[ram_w32_l512_id1_1_addr] <= ram_w32_l512_id1_1_wdata;
        ram_w32_l512_id1_1_rdata_out <= ram_w32_l512_id1_1_wdata;
      end else begin
        ram_w32_l512_id1_1_rdata_out <= mem[ram_w32_l512_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id2
(
  input CLK,
  input [9-1:0] ram_w32_l512_id2_0_addr,
  output [32-1:0] ram_w32_l512_id2_0_rdata,
  input [32-1:0] ram_w32_l512_id2_0_wdata,
  input ram_w32_l512_id2_0_wenable,
  input ram_w32_l512_id2_0_enable,
  input [9-1:0] ram_w32_l512_id2_1_addr,
  output [32-1:0] ram_w32_l512_id2_1_rdata,
  input [32-1:0] ram_w32_l512_id2_1_wdata,
  input ram_w32_l512_id2_1_wenable,
  input ram_w32_l512_id2_1_enable
);

  reg [32-1:0] ram_w32_l512_id2_0_rdata_out;
  assign ram_w32_l512_id2_0_rdata = ram_w32_l512_id2_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id2_1_rdata_out;
  assign ram_w32_l512_id2_1_rdata = ram_w32_l512_id2_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id2_0_enable) begin
      if(ram_w32_l512_id2_0_wenable) begin
        mem[ram_w32_l512_id2_0_addr] <= ram_w32_l512_id2_0_wdata;
        ram_w32_l512_id2_0_rdata_out <= ram_w32_l512_id2_0_wdata;
      end else begin
        ram_w32_l512_id2_0_rdata_out <= mem[ram_w32_l512_id2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id2_1_enable) begin
      if(ram_w32_l512_id2_1_wenable) begin
        mem[ram_w32_l512_id2_1_addr] <= ram_w32_l512_id2_1_wdata;
        ram_w32_l512_id2_1_rdata_out <= ram_w32_l512_id2_1_wdata;
      end else begin
        ram_w32_l512_id2_1_rdata_out <= mem[ram_w32_l512_id2_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id3
(
  input CLK,
  input [9-1:0] ram_w32_l512_id3_0_addr,
  output [32-1:0] ram_w32_l512_id3_0_rdata,
  input [32-1:0] ram_w32_l512_id3_0_wdata,
  input ram_w32_l512_id3_0_wenable,
  input ram_w32_l512_id3_0_enable,
  input [9-1:0] ram_w32_l512_id3_1_addr,
  output [32-1:0] ram_w32_l512_id3_1_rdata,
  input [32-1:0] ram_w32_l512_id3_1_wdata,
  input ram_w32_l512_id3_1_wenable,
  input ram_w32_l512_id3_1_enable
);

  reg [32-1:0] ram_w32_l512_id3_0_rdata_out;
  assign ram_w32_l512_id3_0_rdata = ram_w32_l512_id3_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id3_1_rdata_out;
  assign ram_w32_l512_id3_1_rdata = ram_w32_l512_id3_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id3_0_enable) begin
      if(ram_w32_l512_id3_0_wenable) begin
        mem[ram_w32_l512_id3_0_addr] <= ram_w32_l512_id3_0_wdata;
        ram_w32_l512_id3_0_rdata_out <= ram_w32_l512_id3_0_wdata;
      end else begin
        ram_w32_l512_id3_0_rdata_out <= mem[ram_w32_l512_id3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id3_1_enable) begin
      if(ram_w32_l512_id3_1_wenable) begin
        mem[ram_w32_l512_id3_1_addr] <= ram_w32_l512_id3_1_wdata;
        ram_w32_l512_id3_1_rdata_out <= ram_w32_l512_id3_1_wdata;
      end else begin
        ram_w32_l512_id3_1_rdata_out <= mem[ram_w32_l512_id3_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id4
(
  input CLK,
  input [9-1:0] ram_w32_l512_id4_0_addr,
  output [32-1:0] ram_w32_l512_id4_0_rdata,
  input [32-1:0] ram_w32_l512_id4_0_wdata,
  input ram_w32_l512_id4_0_wenable,
  input ram_w32_l512_id4_0_enable,
  input [9-1:0] ram_w32_l512_id4_1_addr,
  output [32-1:0] ram_w32_l512_id4_1_rdata,
  input [32-1:0] ram_w32_l512_id4_1_wdata,
  input ram_w32_l512_id4_1_wenable,
  input ram_w32_l512_id4_1_enable
);

  reg [32-1:0] ram_w32_l512_id4_0_rdata_out;
  assign ram_w32_l512_id4_0_rdata = ram_w32_l512_id4_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id4_1_rdata_out;
  assign ram_w32_l512_id4_1_rdata = ram_w32_l512_id4_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id4_0_enable) begin
      if(ram_w32_l512_id4_0_wenable) begin
        mem[ram_w32_l512_id4_0_addr] <= ram_w32_l512_id4_0_wdata;
        ram_w32_l512_id4_0_rdata_out <= ram_w32_l512_id4_0_wdata;
      end else begin
        ram_w32_l512_id4_0_rdata_out <= mem[ram_w32_l512_id4_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id4_1_enable) begin
      if(ram_w32_l512_id4_1_wenable) begin
        mem[ram_w32_l512_id4_1_addr] <= ram_w32_l512_id4_1_wdata;
        ram_w32_l512_id4_1_rdata_out <= ram_w32_l512_id4_1_wdata;
      end else begin
        ram_w32_l512_id4_1_rdata_out <= mem[ram_w32_l512_id4_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id5
(
  input CLK,
  input [9-1:0] ram_w32_l512_id5_0_addr,
  output [32-1:0] ram_w32_l512_id5_0_rdata,
  input [32-1:0] ram_w32_l512_id5_0_wdata,
  input ram_w32_l512_id5_0_wenable,
  input ram_w32_l512_id5_0_enable,
  input [9-1:0] ram_w32_l512_id5_1_addr,
  output [32-1:0] ram_w32_l512_id5_1_rdata,
  input [32-1:0] ram_w32_l512_id5_1_wdata,
  input ram_w32_l512_id5_1_wenable,
  input ram_w32_l512_id5_1_enable
);

  reg [32-1:0] ram_w32_l512_id5_0_rdata_out;
  assign ram_w32_l512_id5_0_rdata = ram_w32_l512_id5_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id5_1_rdata_out;
  assign ram_w32_l512_id5_1_rdata = ram_w32_l512_id5_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id5_0_enable) begin
      if(ram_w32_l512_id5_0_wenable) begin
        mem[ram_w32_l512_id5_0_addr] <= ram_w32_l512_id5_0_wdata;
        ram_w32_l512_id5_0_rdata_out <= ram_w32_l512_id5_0_wdata;
      end else begin
        ram_w32_l512_id5_0_rdata_out <= mem[ram_w32_l512_id5_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id5_1_enable) begin
      if(ram_w32_l512_id5_1_wenable) begin
        mem[ram_w32_l512_id5_1_addr] <= ram_w32_l512_id5_1_wdata;
        ram_w32_l512_id5_1_rdata_out <= ram_w32_l512_id5_1_wdata;
      end else begin
        ram_w32_l512_id5_1_rdata_out <= mem[ram_w32_l512_id5_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id6
(
  input CLK,
  input [9-1:0] ram_w32_l512_id6_0_addr,
  output [32-1:0] ram_w32_l512_id6_0_rdata,
  input [32-1:0] ram_w32_l512_id6_0_wdata,
  input ram_w32_l512_id6_0_wenable,
  input ram_w32_l512_id6_0_enable,
  input [9-1:0] ram_w32_l512_id6_1_addr,
  output [32-1:0] ram_w32_l512_id6_1_rdata,
  input [32-1:0] ram_w32_l512_id6_1_wdata,
  input ram_w32_l512_id6_1_wenable,
  input ram_w32_l512_id6_1_enable
);

  reg [32-1:0] ram_w32_l512_id6_0_rdata_out;
  assign ram_w32_l512_id6_0_rdata = ram_w32_l512_id6_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id6_1_rdata_out;
  assign ram_w32_l512_id6_1_rdata = ram_w32_l512_id6_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id6_0_enable) begin
      if(ram_w32_l512_id6_0_wenable) begin
        mem[ram_w32_l512_id6_0_addr] <= ram_w32_l512_id6_0_wdata;
        ram_w32_l512_id6_0_rdata_out <= ram_w32_l512_id6_0_wdata;
      end else begin
        ram_w32_l512_id6_0_rdata_out <= mem[ram_w32_l512_id6_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id6_1_enable) begin
      if(ram_w32_l512_id6_1_wenable) begin
        mem[ram_w32_l512_id6_1_addr] <= ram_w32_l512_id6_1_wdata;
        ram_w32_l512_id6_1_rdata_out <= ram_w32_l512_id6_1_wdata;
      end else begin
        ram_w32_l512_id6_1_rdata_out <= mem[ram_w32_l512_id6_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id7
(
  input CLK,
  input [9-1:0] ram_w32_l512_id7_0_addr,
  output [32-1:0] ram_w32_l512_id7_0_rdata,
  input [32-1:0] ram_w32_l512_id7_0_wdata,
  input ram_w32_l512_id7_0_wenable,
  input ram_w32_l512_id7_0_enable,
  input [9-1:0] ram_w32_l512_id7_1_addr,
  output [32-1:0] ram_w32_l512_id7_1_rdata,
  input [32-1:0] ram_w32_l512_id7_1_wdata,
  input ram_w32_l512_id7_1_wenable,
  input ram_w32_l512_id7_1_enable
);

  reg [32-1:0] ram_w32_l512_id7_0_rdata_out;
  assign ram_w32_l512_id7_0_rdata = ram_w32_l512_id7_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id7_1_rdata_out;
  assign ram_w32_l512_id7_1_rdata = ram_w32_l512_id7_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id7_0_enable) begin
      if(ram_w32_l512_id7_0_wenable) begin
        mem[ram_w32_l512_id7_0_addr] <= ram_w32_l512_id7_0_wdata;
        ram_w32_l512_id7_0_rdata_out <= ram_w32_l512_id7_0_wdata;
      end else begin
        ram_w32_l512_id7_0_rdata_out <= mem[ram_w32_l512_id7_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id7_1_enable) begin
      if(ram_w32_l512_id7_1_wenable) begin
        mem[ram_w32_l512_id7_1_addr] <= ram_w32_l512_id7_1_wdata;
        ram_w32_l512_id7_1_rdata_out <= ram_w32_l512_id7_1_wdata;
      end else begin
        ram_w32_l512_id7_1_rdata_out <= mem[ram_w32_l512_id7_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l512_id8
(
  input CLK,
  input [9-1:0] ram_w32_l512_id8_0_addr,
  output [32-1:0] ram_w32_l512_id8_0_rdata,
  input [32-1:0] ram_w32_l512_id8_0_wdata,
  input ram_w32_l512_id8_0_wenable,
  input ram_w32_l512_id8_0_enable,
  input [9-1:0] ram_w32_l512_id8_1_addr,
  output [32-1:0] ram_w32_l512_id8_1_rdata,
  input [32-1:0] ram_w32_l512_id8_1_wdata,
  input ram_w32_l512_id8_1_wenable,
  input ram_w32_l512_id8_1_enable
);

  reg [32-1:0] ram_w32_l512_id8_0_rdata_out;
  assign ram_w32_l512_id8_0_rdata = ram_w32_l512_id8_0_rdata_out;
  reg [32-1:0] ram_w32_l512_id8_1_rdata_out;
  assign ram_w32_l512_id8_1_rdata = ram_w32_l512_id8_1_rdata_out;
  reg [32-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w32_l512_id8_0_enable) begin
      if(ram_w32_l512_id8_0_wenable) begin
        mem[ram_w32_l512_id8_0_addr] <= ram_w32_l512_id8_0_wdata;
        ram_w32_l512_id8_0_rdata_out <= ram_w32_l512_id8_0_wdata;
      end else begin
        ram_w32_l512_id8_0_rdata_out <= mem[ram_w32_l512_id8_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l512_id8_1_enable) begin
      if(ram_w32_l512_id8_1_wenable) begin
        mem[ram_w32_l512_id8_1_addr] <= ram_w32_l512_id8_1_wdata;
        ram_w32_l512_id8_1_rdata_out <= ram_w32_l512_id8_1_wdata;
      end else begin
        ram_w32_l512_id8_1_rdata_out <= mem[ram_w32_l512_id8_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l256_id0
(
  input CLK,
  input [8-1:0] ram_w32_l256_id0_0_addr,
  output [32-1:0] ram_w32_l256_id0_0_rdata,
  input [32-1:0] ram_w32_l256_id0_0_wdata,
  input ram_w32_l256_id0_0_wenable,
  input ram_w32_l256_id0_0_enable,
  input [8-1:0] ram_w32_l256_id0_1_addr,
  output [32-1:0] ram_w32_l256_id0_1_rdata,
  input [32-1:0] ram_w32_l256_id0_1_wdata,
  input ram_w32_l256_id0_1_wenable,
  input ram_w32_l256_id0_1_enable
);

  reg [32-1:0] ram_w32_l256_id0_0_rdata_out;
  assign ram_w32_l256_id0_0_rdata = ram_w32_l256_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l256_id0_1_rdata_out;
  assign ram_w32_l256_id0_1_rdata = ram_w32_l256_id0_1_rdata_out;
  reg [32-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w32_l256_id0_0_enable) begin
      if(ram_w32_l256_id0_0_wenable) begin
        mem[ram_w32_l256_id0_0_addr] <= ram_w32_l256_id0_0_wdata;
        ram_w32_l256_id0_0_rdata_out <= ram_w32_l256_id0_0_wdata;
      end else begin
        ram_w32_l256_id0_0_rdata_out <= mem[ram_w32_l256_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l256_id0_1_enable) begin
      if(ram_w32_l256_id0_1_wenable) begin
        mem[ram_w32_l256_id0_1_addr] <= ram_w32_l256_id0_1_wdata;
        ram_w32_l256_id0_1_rdata_out <= ram_w32_l256_id0_1_wdata;
      end else begin
        ram_w32_l256_id0_1_rdata_out <= mem[ram_w32_l256_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l256_id1
(
  input CLK,
  input [8-1:0] ram_w32_l256_id1_0_addr,
  output [32-1:0] ram_w32_l256_id1_0_rdata,
  input [32-1:0] ram_w32_l256_id1_0_wdata,
  input ram_w32_l256_id1_0_wenable,
  input ram_w32_l256_id1_0_enable,
  input [8-1:0] ram_w32_l256_id1_1_addr,
  output [32-1:0] ram_w32_l256_id1_1_rdata,
  input [32-1:0] ram_w32_l256_id1_1_wdata,
  input ram_w32_l256_id1_1_wenable,
  input ram_w32_l256_id1_1_enable
);

  reg [32-1:0] ram_w32_l256_id1_0_rdata_out;
  assign ram_w32_l256_id1_0_rdata = ram_w32_l256_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l256_id1_1_rdata_out;
  assign ram_w32_l256_id1_1_rdata = ram_w32_l256_id1_1_rdata_out;
  reg [32-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w32_l256_id1_0_enable) begin
      if(ram_w32_l256_id1_0_wenable) begin
        mem[ram_w32_l256_id1_0_addr] <= ram_w32_l256_id1_0_wdata;
        ram_w32_l256_id1_0_rdata_out <= ram_w32_l256_id1_0_wdata;
      end else begin
        ram_w32_l256_id1_0_rdata_out <= mem[ram_w32_l256_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l256_id1_1_enable) begin
      if(ram_w32_l256_id1_1_wenable) begin
        mem[ram_w32_l256_id1_1_addr] <= ram_w32_l256_id1_1_wdata;
        ram_w32_l256_id1_1_rdata_out <= ram_w32_l256_id1_1_wdata;
      end else begin
        ram_w32_l256_id1_1_rdata_out <= mem[ram_w32_l256_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id0
(
  input CLK,
  input [7-1:0] ram_w32_l128_id0_0_addr,
  output [32-1:0] ram_w32_l128_id0_0_rdata,
  input [32-1:0] ram_w32_l128_id0_0_wdata,
  input ram_w32_l128_id0_0_wenable,
  input ram_w32_l128_id0_0_enable,
  input [7-1:0] ram_w32_l128_id0_1_addr,
  output [32-1:0] ram_w32_l128_id0_1_rdata,
  input [32-1:0] ram_w32_l128_id0_1_wdata,
  input ram_w32_l128_id0_1_wenable,
  input ram_w32_l128_id0_1_enable
);

  reg [32-1:0] ram_w32_l128_id0_0_rdata_out;
  assign ram_w32_l128_id0_0_rdata = ram_w32_l128_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id0_1_rdata_out;
  assign ram_w32_l128_id0_1_rdata = ram_w32_l128_id0_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id0_0_enable) begin
      if(ram_w32_l128_id0_0_wenable) begin
        mem[ram_w32_l128_id0_0_addr] <= ram_w32_l128_id0_0_wdata;
        ram_w32_l128_id0_0_rdata_out <= ram_w32_l128_id0_0_wdata;
      end else begin
        ram_w32_l128_id0_0_rdata_out <= mem[ram_w32_l128_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id0_1_enable) begin
      if(ram_w32_l128_id0_1_wenable) begin
        mem[ram_w32_l128_id0_1_addr] <= ram_w32_l128_id0_1_wdata;
        ram_w32_l128_id0_1_rdata_out <= ram_w32_l128_id0_1_wdata;
      end else begin
        ram_w32_l128_id0_1_rdata_out <= mem[ram_w32_l128_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id1
(
  input CLK,
  input [7-1:0] ram_w32_l128_id1_0_addr,
  output [32-1:0] ram_w32_l128_id1_0_rdata,
  input [32-1:0] ram_w32_l128_id1_0_wdata,
  input ram_w32_l128_id1_0_wenable,
  input ram_w32_l128_id1_0_enable,
  input [7-1:0] ram_w32_l128_id1_1_addr,
  output [32-1:0] ram_w32_l128_id1_1_rdata,
  input [32-1:0] ram_w32_l128_id1_1_wdata,
  input ram_w32_l128_id1_1_wenable,
  input ram_w32_l128_id1_1_enable
);

  reg [32-1:0] ram_w32_l128_id1_0_rdata_out;
  assign ram_w32_l128_id1_0_rdata = ram_w32_l128_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id1_1_rdata_out;
  assign ram_w32_l128_id1_1_rdata = ram_w32_l128_id1_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id1_0_enable) begin
      if(ram_w32_l128_id1_0_wenable) begin
        mem[ram_w32_l128_id1_0_addr] <= ram_w32_l128_id1_0_wdata;
        ram_w32_l128_id1_0_rdata_out <= ram_w32_l128_id1_0_wdata;
      end else begin
        ram_w32_l128_id1_0_rdata_out <= mem[ram_w32_l128_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id1_1_enable) begin
      if(ram_w32_l128_id1_1_wenable) begin
        mem[ram_w32_l128_id1_1_addr] <= ram_w32_l128_id1_1_wdata;
        ram_w32_l128_id1_1_rdata_out <= ram_w32_l128_id1_1_wdata;
      end else begin
        ram_w32_l128_id1_1_rdata_out <= mem[ram_w32_l128_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id2
(
  input CLK,
  input [7-1:0] ram_w32_l128_id2_0_addr,
  output [32-1:0] ram_w32_l128_id2_0_rdata,
  input [32-1:0] ram_w32_l128_id2_0_wdata,
  input ram_w32_l128_id2_0_wenable,
  input ram_w32_l128_id2_0_enable,
  input [7-1:0] ram_w32_l128_id2_1_addr,
  output [32-1:0] ram_w32_l128_id2_1_rdata,
  input [32-1:0] ram_w32_l128_id2_1_wdata,
  input ram_w32_l128_id2_1_wenable,
  input ram_w32_l128_id2_1_enable
);

  reg [32-1:0] ram_w32_l128_id2_0_rdata_out;
  assign ram_w32_l128_id2_0_rdata = ram_w32_l128_id2_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id2_1_rdata_out;
  assign ram_w32_l128_id2_1_rdata = ram_w32_l128_id2_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id2_0_enable) begin
      if(ram_w32_l128_id2_0_wenable) begin
        mem[ram_w32_l128_id2_0_addr] <= ram_w32_l128_id2_0_wdata;
        ram_w32_l128_id2_0_rdata_out <= ram_w32_l128_id2_0_wdata;
      end else begin
        ram_w32_l128_id2_0_rdata_out <= mem[ram_w32_l128_id2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id2_1_enable) begin
      if(ram_w32_l128_id2_1_wenable) begin
        mem[ram_w32_l128_id2_1_addr] <= ram_w32_l128_id2_1_wdata;
        ram_w32_l128_id2_1_rdata_out <= ram_w32_l128_id2_1_wdata;
      end else begin
        ram_w32_l128_id2_1_rdata_out <= mem[ram_w32_l128_id2_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id3
(
  input CLK,
  input [7-1:0] ram_w32_l128_id3_0_addr,
  output [32-1:0] ram_w32_l128_id3_0_rdata,
  input [32-1:0] ram_w32_l128_id3_0_wdata,
  input ram_w32_l128_id3_0_wenable,
  input ram_w32_l128_id3_0_enable,
  input [7-1:0] ram_w32_l128_id3_1_addr,
  output [32-1:0] ram_w32_l128_id3_1_rdata,
  input [32-1:0] ram_w32_l128_id3_1_wdata,
  input ram_w32_l128_id3_1_wenable,
  input ram_w32_l128_id3_1_enable
);

  reg [32-1:0] ram_w32_l128_id3_0_rdata_out;
  assign ram_w32_l128_id3_0_rdata = ram_w32_l128_id3_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id3_1_rdata_out;
  assign ram_w32_l128_id3_1_rdata = ram_w32_l128_id3_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id3_0_enable) begin
      if(ram_w32_l128_id3_0_wenable) begin
        mem[ram_w32_l128_id3_0_addr] <= ram_w32_l128_id3_0_wdata;
        ram_w32_l128_id3_0_rdata_out <= ram_w32_l128_id3_0_wdata;
      end else begin
        ram_w32_l128_id3_0_rdata_out <= mem[ram_w32_l128_id3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id3_1_enable) begin
      if(ram_w32_l128_id3_1_wenable) begin
        mem[ram_w32_l128_id3_1_addr] <= ram_w32_l128_id3_1_wdata;
        ram_w32_l128_id3_1_rdata_out <= ram_w32_l128_id3_1_wdata;
      end else begin
        ram_w32_l128_id3_1_rdata_out <= mem[ram_w32_l128_id3_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id4
(
  input CLK,
  input [7-1:0] ram_w32_l128_id4_0_addr,
  output [32-1:0] ram_w32_l128_id4_0_rdata,
  input [32-1:0] ram_w32_l128_id4_0_wdata,
  input ram_w32_l128_id4_0_wenable,
  input ram_w32_l128_id4_0_enable,
  input [7-1:0] ram_w32_l128_id4_1_addr,
  output [32-1:0] ram_w32_l128_id4_1_rdata,
  input [32-1:0] ram_w32_l128_id4_1_wdata,
  input ram_w32_l128_id4_1_wenable,
  input ram_w32_l128_id4_1_enable
);

  reg [32-1:0] ram_w32_l128_id4_0_rdata_out;
  assign ram_w32_l128_id4_0_rdata = ram_w32_l128_id4_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id4_1_rdata_out;
  assign ram_w32_l128_id4_1_rdata = ram_w32_l128_id4_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id4_0_enable) begin
      if(ram_w32_l128_id4_0_wenable) begin
        mem[ram_w32_l128_id4_0_addr] <= ram_w32_l128_id4_0_wdata;
        ram_w32_l128_id4_0_rdata_out <= ram_w32_l128_id4_0_wdata;
      end else begin
        ram_w32_l128_id4_0_rdata_out <= mem[ram_w32_l128_id4_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id4_1_enable) begin
      if(ram_w32_l128_id4_1_wenable) begin
        mem[ram_w32_l128_id4_1_addr] <= ram_w32_l128_id4_1_wdata;
        ram_w32_l128_id4_1_rdata_out <= ram_w32_l128_id4_1_wdata;
      end else begin
        ram_w32_l128_id4_1_rdata_out <= mem[ram_w32_l128_id4_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id5
(
  input CLK,
  input [7-1:0] ram_w32_l128_id5_0_addr,
  output [32-1:0] ram_w32_l128_id5_0_rdata,
  input [32-1:0] ram_w32_l128_id5_0_wdata,
  input ram_w32_l128_id5_0_wenable,
  input ram_w32_l128_id5_0_enable,
  input [7-1:0] ram_w32_l128_id5_1_addr,
  output [32-1:0] ram_w32_l128_id5_1_rdata,
  input [32-1:0] ram_w32_l128_id5_1_wdata,
  input ram_w32_l128_id5_1_wenable,
  input ram_w32_l128_id5_1_enable
);

  reg [32-1:0] ram_w32_l128_id5_0_rdata_out;
  assign ram_w32_l128_id5_0_rdata = ram_w32_l128_id5_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id5_1_rdata_out;
  assign ram_w32_l128_id5_1_rdata = ram_w32_l128_id5_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id5_0_enable) begin
      if(ram_w32_l128_id5_0_wenable) begin
        mem[ram_w32_l128_id5_0_addr] <= ram_w32_l128_id5_0_wdata;
        ram_w32_l128_id5_0_rdata_out <= ram_w32_l128_id5_0_wdata;
      end else begin
        ram_w32_l128_id5_0_rdata_out <= mem[ram_w32_l128_id5_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id5_1_enable) begin
      if(ram_w32_l128_id5_1_wenable) begin
        mem[ram_w32_l128_id5_1_addr] <= ram_w32_l128_id5_1_wdata;
        ram_w32_l128_id5_1_rdata_out <= ram_w32_l128_id5_1_wdata;
      end else begin
        ram_w32_l128_id5_1_rdata_out <= mem[ram_w32_l128_id5_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id6
(
  input CLK,
  input [7-1:0] ram_w32_l128_id6_0_addr,
  output [32-1:0] ram_w32_l128_id6_0_rdata,
  input [32-1:0] ram_w32_l128_id6_0_wdata,
  input ram_w32_l128_id6_0_wenable,
  input ram_w32_l128_id6_0_enable,
  input [7-1:0] ram_w32_l128_id6_1_addr,
  output [32-1:0] ram_w32_l128_id6_1_rdata,
  input [32-1:0] ram_w32_l128_id6_1_wdata,
  input ram_w32_l128_id6_1_wenable,
  input ram_w32_l128_id6_1_enable
);

  reg [32-1:0] ram_w32_l128_id6_0_rdata_out;
  assign ram_w32_l128_id6_0_rdata = ram_w32_l128_id6_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id6_1_rdata_out;
  assign ram_w32_l128_id6_1_rdata = ram_w32_l128_id6_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id6_0_enable) begin
      if(ram_w32_l128_id6_0_wenable) begin
        mem[ram_w32_l128_id6_0_addr] <= ram_w32_l128_id6_0_wdata;
        ram_w32_l128_id6_0_rdata_out <= ram_w32_l128_id6_0_wdata;
      end else begin
        ram_w32_l128_id6_0_rdata_out <= mem[ram_w32_l128_id6_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id6_1_enable) begin
      if(ram_w32_l128_id6_1_wenable) begin
        mem[ram_w32_l128_id6_1_addr] <= ram_w32_l128_id6_1_wdata;
        ram_w32_l128_id6_1_rdata_out <= ram_w32_l128_id6_1_wdata;
      end else begin
        ram_w32_l128_id6_1_rdata_out <= mem[ram_w32_l128_id6_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id7
(
  input CLK,
  input [7-1:0] ram_w32_l128_id7_0_addr,
  output [32-1:0] ram_w32_l128_id7_0_rdata,
  input [32-1:0] ram_w32_l128_id7_0_wdata,
  input ram_w32_l128_id7_0_wenable,
  input ram_w32_l128_id7_0_enable,
  input [7-1:0] ram_w32_l128_id7_1_addr,
  output [32-1:0] ram_w32_l128_id7_1_rdata,
  input [32-1:0] ram_w32_l128_id7_1_wdata,
  input ram_w32_l128_id7_1_wenable,
  input ram_w32_l128_id7_1_enable
);

  reg [32-1:0] ram_w32_l128_id7_0_rdata_out;
  assign ram_w32_l128_id7_0_rdata = ram_w32_l128_id7_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id7_1_rdata_out;
  assign ram_w32_l128_id7_1_rdata = ram_w32_l128_id7_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id7_0_enable) begin
      if(ram_w32_l128_id7_0_wenable) begin
        mem[ram_w32_l128_id7_0_addr] <= ram_w32_l128_id7_0_wdata;
        ram_w32_l128_id7_0_rdata_out <= ram_w32_l128_id7_0_wdata;
      end else begin
        ram_w32_l128_id7_0_rdata_out <= mem[ram_w32_l128_id7_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id7_1_enable) begin
      if(ram_w32_l128_id7_1_wenable) begin
        mem[ram_w32_l128_id7_1_addr] <= ram_w32_l128_id7_1_wdata;
        ram_w32_l128_id7_1_rdata_out <= ram_w32_l128_id7_1_wdata;
      end else begin
        ram_w32_l128_id7_1_rdata_out <= mem[ram_w32_l128_id7_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id8
(
  input CLK,
  input [7-1:0] ram_w32_l128_id8_0_addr,
  output [32-1:0] ram_w32_l128_id8_0_rdata,
  input [32-1:0] ram_w32_l128_id8_0_wdata,
  input ram_w32_l128_id8_0_wenable,
  input ram_w32_l128_id8_0_enable,
  input [7-1:0] ram_w32_l128_id8_1_addr,
  output [32-1:0] ram_w32_l128_id8_1_rdata,
  input [32-1:0] ram_w32_l128_id8_1_wdata,
  input ram_w32_l128_id8_1_wenable,
  input ram_w32_l128_id8_1_enable
);

  reg [32-1:0] ram_w32_l128_id8_0_rdata_out;
  assign ram_w32_l128_id8_0_rdata = ram_w32_l128_id8_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id8_1_rdata_out;
  assign ram_w32_l128_id8_1_rdata = ram_w32_l128_id8_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id8_0_enable) begin
      if(ram_w32_l128_id8_0_wenable) begin
        mem[ram_w32_l128_id8_0_addr] <= ram_w32_l128_id8_0_wdata;
        ram_w32_l128_id8_0_rdata_out <= ram_w32_l128_id8_0_wdata;
      end else begin
        ram_w32_l128_id8_0_rdata_out <= mem[ram_w32_l128_id8_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id8_1_enable) begin
      if(ram_w32_l128_id8_1_wenable) begin
        mem[ram_w32_l128_id8_1_addr] <= ram_w32_l128_id8_1_wdata;
        ram_w32_l128_id8_1_rdata_out <= ram_w32_l128_id8_1_wdata;
      end else begin
        ram_w32_l128_id8_1_rdata_out <= mem[ram_w32_l128_id8_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id9
(
  input CLK,
  input [7-1:0] ram_w32_l128_id9_0_addr,
  output [32-1:0] ram_w32_l128_id9_0_rdata,
  input [32-1:0] ram_w32_l128_id9_0_wdata,
  input ram_w32_l128_id9_0_wenable,
  input ram_w32_l128_id9_0_enable,
  input [7-1:0] ram_w32_l128_id9_1_addr,
  output [32-1:0] ram_w32_l128_id9_1_rdata,
  input [32-1:0] ram_w32_l128_id9_1_wdata,
  input ram_w32_l128_id9_1_wenable,
  input ram_w32_l128_id9_1_enable
);

  reg [32-1:0] ram_w32_l128_id9_0_rdata_out;
  assign ram_w32_l128_id9_0_rdata = ram_w32_l128_id9_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id9_1_rdata_out;
  assign ram_w32_l128_id9_1_rdata = ram_w32_l128_id9_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id9_0_enable) begin
      if(ram_w32_l128_id9_0_wenable) begin
        mem[ram_w32_l128_id9_0_addr] <= ram_w32_l128_id9_0_wdata;
        ram_w32_l128_id9_0_rdata_out <= ram_w32_l128_id9_0_wdata;
      end else begin
        ram_w32_l128_id9_0_rdata_out <= mem[ram_w32_l128_id9_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id9_1_enable) begin
      if(ram_w32_l128_id9_1_wenable) begin
        mem[ram_w32_l128_id9_1_addr] <= ram_w32_l128_id9_1_wdata;
        ram_w32_l128_id9_1_rdata_out <= ram_w32_l128_id9_1_wdata;
      end else begin
        ram_w32_l128_id9_1_rdata_out <= mem[ram_w32_l128_id9_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id10
(
  input CLK,
  input [7-1:0] ram_w32_l128_id10_0_addr,
  output [32-1:0] ram_w32_l128_id10_0_rdata,
  input [32-1:0] ram_w32_l128_id10_0_wdata,
  input ram_w32_l128_id10_0_wenable,
  input ram_w32_l128_id10_0_enable,
  input [7-1:0] ram_w32_l128_id10_1_addr,
  output [32-1:0] ram_w32_l128_id10_1_rdata,
  input [32-1:0] ram_w32_l128_id10_1_wdata,
  input ram_w32_l128_id10_1_wenable,
  input ram_w32_l128_id10_1_enable
);

  reg [32-1:0] ram_w32_l128_id10_0_rdata_out;
  assign ram_w32_l128_id10_0_rdata = ram_w32_l128_id10_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id10_1_rdata_out;
  assign ram_w32_l128_id10_1_rdata = ram_w32_l128_id10_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id10_0_enable) begin
      if(ram_w32_l128_id10_0_wenable) begin
        mem[ram_w32_l128_id10_0_addr] <= ram_w32_l128_id10_0_wdata;
        ram_w32_l128_id10_0_rdata_out <= ram_w32_l128_id10_0_wdata;
      end else begin
        ram_w32_l128_id10_0_rdata_out <= mem[ram_w32_l128_id10_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id10_1_enable) begin
      if(ram_w32_l128_id10_1_wenable) begin
        mem[ram_w32_l128_id10_1_addr] <= ram_w32_l128_id10_1_wdata;
        ram_w32_l128_id10_1_rdata_out <= ram_w32_l128_id10_1_wdata;
      end else begin
        ram_w32_l128_id10_1_rdata_out <= mem[ram_w32_l128_id10_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id11
(
  input CLK,
  input [7-1:0] ram_w32_l128_id11_0_addr,
  output [32-1:0] ram_w32_l128_id11_0_rdata,
  input [32-1:0] ram_w32_l128_id11_0_wdata,
  input ram_w32_l128_id11_0_wenable,
  input ram_w32_l128_id11_0_enable,
  input [7-1:0] ram_w32_l128_id11_1_addr,
  output [32-1:0] ram_w32_l128_id11_1_rdata,
  input [32-1:0] ram_w32_l128_id11_1_wdata,
  input ram_w32_l128_id11_1_wenable,
  input ram_w32_l128_id11_1_enable
);

  reg [32-1:0] ram_w32_l128_id11_0_rdata_out;
  assign ram_w32_l128_id11_0_rdata = ram_w32_l128_id11_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id11_1_rdata_out;
  assign ram_w32_l128_id11_1_rdata = ram_w32_l128_id11_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id11_0_enable) begin
      if(ram_w32_l128_id11_0_wenable) begin
        mem[ram_w32_l128_id11_0_addr] <= ram_w32_l128_id11_0_wdata;
        ram_w32_l128_id11_0_rdata_out <= ram_w32_l128_id11_0_wdata;
      end else begin
        ram_w32_l128_id11_0_rdata_out <= mem[ram_w32_l128_id11_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id11_1_enable) begin
      if(ram_w32_l128_id11_1_wenable) begin
        mem[ram_w32_l128_id11_1_addr] <= ram_w32_l128_id11_1_wdata;
        ram_w32_l128_id11_1_rdata_out <= ram_w32_l128_id11_1_wdata;
      end else begin
        ram_w32_l128_id11_1_rdata_out <= mem[ram_w32_l128_id11_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id12
(
  input CLK,
  input [7-1:0] ram_w32_l128_id12_0_addr,
  output [32-1:0] ram_w32_l128_id12_0_rdata,
  input [32-1:0] ram_w32_l128_id12_0_wdata,
  input ram_w32_l128_id12_0_wenable,
  input ram_w32_l128_id12_0_enable,
  input [7-1:0] ram_w32_l128_id12_1_addr,
  output [32-1:0] ram_w32_l128_id12_1_rdata,
  input [32-1:0] ram_w32_l128_id12_1_wdata,
  input ram_w32_l128_id12_1_wenable,
  input ram_w32_l128_id12_1_enable
);

  reg [32-1:0] ram_w32_l128_id12_0_rdata_out;
  assign ram_w32_l128_id12_0_rdata = ram_w32_l128_id12_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id12_1_rdata_out;
  assign ram_w32_l128_id12_1_rdata = ram_w32_l128_id12_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id12_0_enable) begin
      if(ram_w32_l128_id12_0_wenable) begin
        mem[ram_w32_l128_id12_0_addr] <= ram_w32_l128_id12_0_wdata;
        ram_w32_l128_id12_0_rdata_out <= ram_w32_l128_id12_0_wdata;
      end else begin
        ram_w32_l128_id12_0_rdata_out <= mem[ram_w32_l128_id12_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id12_1_enable) begin
      if(ram_w32_l128_id12_1_wenable) begin
        mem[ram_w32_l128_id12_1_addr] <= ram_w32_l128_id12_1_wdata;
        ram_w32_l128_id12_1_rdata_out <= ram_w32_l128_id12_1_wdata;
      end else begin
        ram_w32_l128_id12_1_rdata_out <= mem[ram_w32_l128_id12_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id13
(
  input CLK,
  input [7-1:0] ram_w32_l128_id13_0_addr,
  output [32-1:0] ram_w32_l128_id13_0_rdata,
  input [32-1:0] ram_w32_l128_id13_0_wdata,
  input ram_w32_l128_id13_0_wenable,
  input ram_w32_l128_id13_0_enable,
  input [7-1:0] ram_w32_l128_id13_1_addr,
  output [32-1:0] ram_w32_l128_id13_1_rdata,
  input [32-1:0] ram_w32_l128_id13_1_wdata,
  input ram_w32_l128_id13_1_wenable,
  input ram_w32_l128_id13_1_enable
);

  reg [32-1:0] ram_w32_l128_id13_0_rdata_out;
  assign ram_w32_l128_id13_0_rdata = ram_w32_l128_id13_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id13_1_rdata_out;
  assign ram_w32_l128_id13_1_rdata = ram_w32_l128_id13_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id13_0_enable) begin
      if(ram_w32_l128_id13_0_wenable) begin
        mem[ram_w32_l128_id13_0_addr] <= ram_w32_l128_id13_0_wdata;
        ram_w32_l128_id13_0_rdata_out <= ram_w32_l128_id13_0_wdata;
      end else begin
        ram_w32_l128_id13_0_rdata_out <= mem[ram_w32_l128_id13_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id13_1_enable) begin
      if(ram_w32_l128_id13_1_wenable) begin
        mem[ram_w32_l128_id13_1_addr] <= ram_w32_l128_id13_1_wdata;
        ram_w32_l128_id13_1_rdata_out <= ram_w32_l128_id13_1_wdata;
      end else begin
        ram_w32_l128_id13_1_rdata_out <= mem[ram_w32_l128_id13_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id14
(
  input CLK,
  input [7-1:0] ram_w32_l128_id14_0_addr,
  output [32-1:0] ram_w32_l128_id14_0_rdata,
  input [32-1:0] ram_w32_l128_id14_0_wdata,
  input ram_w32_l128_id14_0_wenable,
  input ram_w32_l128_id14_0_enable,
  input [7-1:0] ram_w32_l128_id14_1_addr,
  output [32-1:0] ram_w32_l128_id14_1_rdata,
  input [32-1:0] ram_w32_l128_id14_1_wdata,
  input ram_w32_l128_id14_1_wenable,
  input ram_w32_l128_id14_1_enable
);

  reg [32-1:0] ram_w32_l128_id14_0_rdata_out;
  assign ram_w32_l128_id14_0_rdata = ram_w32_l128_id14_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id14_1_rdata_out;
  assign ram_w32_l128_id14_1_rdata = ram_w32_l128_id14_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id14_0_enable) begin
      if(ram_w32_l128_id14_0_wenable) begin
        mem[ram_w32_l128_id14_0_addr] <= ram_w32_l128_id14_0_wdata;
        ram_w32_l128_id14_0_rdata_out <= ram_w32_l128_id14_0_wdata;
      end else begin
        ram_w32_l128_id14_0_rdata_out <= mem[ram_w32_l128_id14_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id14_1_enable) begin
      if(ram_w32_l128_id14_1_wenable) begin
        mem[ram_w32_l128_id14_1_addr] <= ram_w32_l128_id14_1_wdata;
        ram_w32_l128_id14_1_rdata_out <= ram_w32_l128_id14_1_wdata;
      end else begin
        ram_w32_l128_id14_1_rdata_out <= mem[ram_w32_l128_id14_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id15
(
  input CLK,
  input [7-1:0] ram_w32_l128_id15_0_addr,
  output [32-1:0] ram_w32_l128_id15_0_rdata,
  input [32-1:0] ram_w32_l128_id15_0_wdata,
  input ram_w32_l128_id15_0_wenable,
  input ram_w32_l128_id15_0_enable,
  input [7-1:0] ram_w32_l128_id15_1_addr,
  output [32-1:0] ram_w32_l128_id15_1_rdata,
  input [32-1:0] ram_w32_l128_id15_1_wdata,
  input ram_w32_l128_id15_1_wenable,
  input ram_w32_l128_id15_1_enable
);

  reg [32-1:0] ram_w32_l128_id15_0_rdata_out;
  assign ram_w32_l128_id15_0_rdata = ram_w32_l128_id15_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id15_1_rdata_out;
  assign ram_w32_l128_id15_1_rdata = ram_w32_l128_id15_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id15_0_enable) begin
      if(ram_w32_l128_id15_0_wenable) begin
        mem[ram_w32_l128_id15_0_addr] <= ram_w32_l128_id15_0_wdata;
        ram_w32_l128_id15_0_rdata_out <= ram_w32_l128_id15_0_wdata;
      end else begin
        ram_w32_l128_id15_0_rdata_out <= mem[ram_w32_l128_id15_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id15_1_enable) begin
      if(ram_w32_l128_id15_1_wenable) begin
        mem[ram_w32_l128_id15_1_addr] <= ram_w32_l128_id15_1_wdata;
        ram_w32_l128_id15_1_rdata_out <= ram_w32_l128_id15_1_wdata;
      end else begin
        ram_w32_l128_id15_1_rdata_out <= mem[ram_w32_l128_id15_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id16
(
  input CLK,
  input [7-1:0] ram_w32_l128_id16_0_addr,
  output [32-1:0] ram_w32_l128_id16_0_rdata,
  input [32-1:0] ram_w32_l128_id16_0_wdata,
  input ram_w32_l128_id16_0_wenable,
  input ram_w32_l128_id16_0_enable,
  input [7-1:0] ram_w32_l128_id16_1_addr,
  output [32-1:0] ram_w32_l128_id16_1_rdata,
  input [32-1:0] ram_w32_l128_id16_1_wdata,
  input ram_w32_l128_id16_1_wenable,
  input ram_w32_l128_id16_1_enable
);

  reg [32-1:0] ram_w32_l128_id16_0_rdata_out;
  assign ram_w32_l128_id16_0_rdata = ram_w32_l128_id16_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id16_1_rdata_out;
  assign ram_w32_l128_id16_1_rdata = ram_w32_l128_id16_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id16_0_enable) begin
      if(ram_w32_l128_id16_0_wenable) begin
        mem[ram_w32_l128_id16_0_addr] <= ram_w32_l128_id16_0_wdata;
        ram_w32_l128_id16_0_rdata_out <= ram_w32_l128_id16_0_wdata;
      end else begin
        ram_w32_l128_id16_0_rdata_out <= mem[ram_w32_l128_id16_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id16_1_enable) begin
      if(ram_w32_l128_id16_1_wenable) begin
        mem[ram_w32_l128_id16_1_addr] <= ram_w32_l128_id16_1_wdata;
        ram_w32_l128_id16_1_rdata_out <= ram_w32_l128_id16_1_wdata;
      end else begin
        ram_w32_l128_id16_1_rdata_out <= mem[ram_w32_l128_id16_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id17
(
  input CLK,
  input [7-1:0] ram_w32_l128_id17_0_addr,
  output [32-1:0] ram_w32_l128_id17_0_rdata,
  input [32-1:0] ram_w32_l128_id17_0_wdata,
  input ram_w32_l128_id17_0_wenable,
  input ram_w32_l128_id17_0_enable,
  input [7-1:0] ram_w32_l128_id17_1_addr,
  output [32-1:0] ram_w32_l128_id17_1_rdata,
  input [32-1:0] ram_w32_l128_id17_1_wdata,
  input ram_w32_l128_id17_1_wenable,
  input ram_w32_l128_id17_1_enable
);

  reg [32-1:0] ram_w32_l128_id17_0_rdata_out;
  assign ram_w32_l128_id17_0_rdata = ram_w32_l128_id17_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id17_1_rdata_out;
  assign ram_w32_l128_id17_1_rdata = ram_w32_l128_id17_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id17_0_enable) begin
      if(ram_w32_l128_id17_0_wenable) begin
        mem[ram_w32_l128_id17_0_addr] <= ram_w32_l128_id17_0_wdata;
        ram_w32_l128_id17_0_rdata_out <= ram_w32_l128_id17_0_wdata;
      end else begin
        ram_w32_l128_id17_0_rdata_out <= mem[ram_w32_l128_id17_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id17_1_enable) begin
      if(ram_w32_l128_id17_1_wenable) begin
        mem[ram_w32_l128_id17_1_addr] <= ram_w32_l128_id17_1_wdata;
        ram_w32_l128_id17_1_rdata_out <= ram_w32_l128_id17_1_wdata;
      end else begin
        ram_w32_l128_id17_1_rdata_out <= mem[ram_w32_l128_id17_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id18
(
  input CLK,
  input [7-1:0] ram_w32_l128_id18_0_addr,
  output [32-1:0] ram_w32_l128_id18_0_rdata,
  input [32-1:0] ram_w32_l128_id18_0_wdata,
  input ram_w32_l128_id18_0_wenable,
  input ram_w32_l128_id18_0_enable,
  input [7-1:0] ram_w32_l128_id18_1_addr,
  output [32-1:0] ram_w32_l128_id18_1_rdata,
  input [32-1:0] ram_w32_l128_id18_1_wdata,
  input ram_w32_l128_id18_1_wenable,
  input ram_w32_l128_id18_1_enable
);

  reg [32-1:0] ram_w32_l128_id18_0_rdata_out;
  assign ram_w32_l128_id18_0_rdata = ram_w32_l128_id18_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id18_1_rdata_out;
  assign ram_w32_l128_id18_1_rdata = ram_w32_l128_id18_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id18_0_enable) begin
      if(ram_w32_l128_id18_0_wenable) begin
        mem[ram_w32_l128_id18_0_addr] <= ram_w32_l128_id18_0_wdata;
        ram_w32_l128_id18_0_rdata_out <= ram_w32_l128_id18_0_wdata;
      end else begin
        ram_w32_l128_id18_0_rdata_out <= mem[ram_w32_l128_id18_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id18_1_enable) begin
      if(ram_w32_l128_id18_1_wenable) begin
        mem[ram_w32_l128_id18_1_addr] <= ram_w32_l128_id18_1_wdata;
        ram_w32_l128_id18_1_rdata_out <= ram_w32_l128_id18_1_wdata;
      end else begin
        ram_w32_l128_id18_1_rdata_out <= mem[ram_w32_l128_id18_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id19
(
  input CLK,
  input [7-1:0] ram_w32_l128_id19_0_addr,
  output [32-1:0] ram_w32_l128_id19_0_rdata,
  input [32-1:0] ram_w32_l128_id19_0_wdata,
  input ram_w32_l128_id19_0_wenable,
  input ram_w32_l128_id19_0_enable,
  input [7-1:0] ram_w32_l128_id19_1_addr,
  output [32-1:0] ram_w32_l128_id19_1_rdata,
  input [32-1:0] ram_w32_l128_id19_1_wdata,
  input ram_w32_l128_id19_1_wenable,
  input ram_w32_l128_id19_1_enable
);

  reg [32-1:0] ram_w32_l128_id19_0_rdata_out;
  assign ram_w32_l128_id19_0_rdata = ram_w32_l128_id19_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id19_1_rdata_out;
  assign ram_w32_l128_id19_1_rdata = ram_w32_l128_id19_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id19_0_enable) begin
      if(ram_w32_l128_id19_0_wenable) begin
        mem[ram_w32_l128_id19_0_addr] <= ram_w32_l128_id19_0_wdata;
        ram_w32_l128_id19_0_rdata_out <= ram_w32_l128_id19_0_wdata;
      end else begin
        ram_w32_l128_id19_0_rdata_out <= mem[ram_w32_l128_id19_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id19_1_enable) begin
      if(ram_w32_l128_id19_1_wenable) begin
        mem[ram_w32_l128_id19_1_addr] <= ram_w32_l128_id19_1_wdata;
        ram_w32_l128_id19_1_rdata_out <= ram_w32_l128_id19_1_wdata;
      end else begin
        ram_w32_l128_id19_1_rdata_out <= mem[ram_w32_l128_id19_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id20
(
  input CLK,
  input [7-1:0] ram_w32_l128_id20_0_addr,
  output [32-1:0] ram_w32_l128_id20_0_rdata,
  input [32-1:0] ram_w32_l128_id20_0_wdata,
  input ram_w32_l128_id20_0_wenable,
  input ram_w32_l128_id20_0_enable,
  input [7-1:0] ram_w32_l128_id20_1_addr,
  output [32-1:0] ram_w32_l128_id20_1_rdata,
  input [32-1:0] ram_w32_l128_id20_1_wdata,
  input ram_w32_l128_id20_1_wenable,
  input ram_w32_l128_id20_1_enable
);

  reg [32-1:0] ram_w32_l128_id20_0_rdata_out;
  assign ram_w32_l128_id20_0_rdata = ram_w32_l128_id20_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id20_1_rdata_out;
  assign ram_w32_l128_id20_1_rdata = ram_w32_l128_id20_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id20_0_enable) begin
      if(ram_w32_l128_id20_0_wenable) begin
        mem[ram_w32_l128_id20_0_addr] <= ram_w32_l128_id20_0_wdata;
        ram_w32_l128_id20_0_rdata_out <= ram_w32_l128_id20_0_wdata;
      end else begin
        ram_w32_l128_id20_0_rdata_out <= mem[ram_w32_l128_id20_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id20_1_enable) begin
      if(ram_w32_l128_id20_1_wenable) begin
        mem[ram_w32_l128_id20_1_addr] <= ram_w32_l128_id20_1_wdata;
        ram_w32_l128_id20_1_rdata_out <= ram_w32_l128_id20_1_wdata;
      end else begin
        ram_w32_l128_id20_1_rdata_out <= mem[ram_w32_l128_id20_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id21
(
  input CLK,
  input [7-1:0] ram_w32_l128_id21_0_addr,
  output [32-1:0] ram_w32_l128_id21_0_rdata,
  input [32-1:0] ram_w32_l128_id21_0_wdata,
  input ram_w32_l128_id21_0_wenable,
  input ram_w32_l128_id21_0_enable,
  input [7-1:0] ram_w32_l128_id21_1_addr,
  output [32-1:0] ram_w32_l128_id21_1_rdata,
  input [32-1:0] ram_w32_l128_id21_1_wdata,
  input ram_w32_l128_id21_1_wenable,
  input ram_w32_l128_id21_1_enable
);

  reg [32-1:0] ram_w32_l128_id21_0_rdata_out;
  assign ram_w32_l128_id21_0_rdata = ram_w32_l128_id21_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id21_1_rdata_out;
  assign ram_w32_l128_id21_1_rdata = ram_w32_l128_id21_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id21_0_enable) begin
      if(ram_w32_l128_id21_0_wenable) begin
        mem[ram_w32_l128_id21_0_addr] <= ram_w32_l128_id21_0_wdata;
        ram_w32_l128_id21_0_rdata_out <= ram_w32_l128_id21_0_wdata;
      end else begin
        ram_w32_l128_id21_0_rdata_out <= mem[ram_w32_l128_id21_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id21_1_enable) begin
      if(ram_w32_l128_id21_1_wenable) begin
        mem[ram_w32_l128_id21_1_addr] <= ram_w32_l128_id21_1_wdata;
        ram_w32_l128_id21_1_rdata_out <= ram_w32_l128_id21_1_wdata;
      end else begin
        ram_w32_l128_id21_1_rdata_out <= mem[ram_w32_l128_id21_1_addr];
      end
    end 
  end


endmodule



module madd_0
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_0
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_0
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_1
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_1
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_1
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_2
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_2
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_2
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_3
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_3
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_3
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_4
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_4
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_4
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_5
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_5
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_5
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_6
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_6
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_6
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_7
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_7
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_7
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_8
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_8
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_8
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_9
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_9
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_9
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_10
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_10
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_10
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_11
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_11
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_11
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_12
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_12
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_12
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_13
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_13
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_13
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_14
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_14
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_14
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_15
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_15
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_15
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_16
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_16
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_16
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_17
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_17
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_17
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_0
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);


  multiplier_core_0
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_0
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);

  reg signed [64-1:0] _a;
  reg signed [16-1:0] _b;
  wire signed [80-1:0] _mul;
  reg signed [80-1:0] _pipe_mul0;
  reg signed [80-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule



module madd_18
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_18
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_18
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_19
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_19
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_19
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_20
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_20
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_20
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_21
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_21
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_21
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_22
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_22
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_22
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_23
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_23
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_23
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_24
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_24
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_24
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_25
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_25
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_25
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_26
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_26
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_26
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_27
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_27
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_27
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_28
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_28
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_28
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_29
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_29
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_29
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_30
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_30
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_30
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_31
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_31
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_31
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_32
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_32
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_32
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_33
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_33
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_33
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_34
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_34
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_34
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_35
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_35
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_35
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_1
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);


  multiplier_core_1
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_1
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);

  reg signed [64-1:0] _a;
  reg signed [16-1:0] _b;
  wire signed [80-1:0] _mul;
  reg signed [80-1:0] _pipe_mul0;
  reg signed [80-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule

